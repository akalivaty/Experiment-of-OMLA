//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n462), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n467), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT65), .A3(G137), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n464), .A2(new_n467), .ZN(new_n479));
  MUX2_X1   g054(.A(G100), .B(G112), .S(G2105), .Z(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G124), .B1(G2104), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(new_n472), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n472), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n475), .A2(new_n488), .A3(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  MUX2_X1   g065(.A(G102), .B(G114), .S(G2105), .Z(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n471), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n479), .A2(G126), .B1(G2104), .B2(new_n491), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n490), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n503), .A2(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT69), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n511), .B2(new_n517), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n502), .A2(G51), .A3(G543), .ZN(new_n521));
  AND3_X1   g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n506), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n502), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  OAI211_X1 g110(.A(G52), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT72), .B(G90), .Z(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n509), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(G64), .B1(new_n506), .B2(new_n505), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n512), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n513), .A2(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n512), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(G43), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n509), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n502), .A2(new_n560), .A3(G53), .A4(G543), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n513), .A2(new_n502), .A3(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n513), .B2(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(new_n512), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n557), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n564), .B1(new_n531), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n505), .ZN(new_n571));
  NAND2_X1  g146(.A1(KEYINPUT5), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(new_n512), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n570), .A2(G651), .B1(new_n576), .B2(G91), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n559), .A2(new_n561), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(KEYINPUT74), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n568), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  NAND2_X1  g159(.A1(new_n576), .A2(G87), .ZN(new_n585));
  INV_X1    g160(.A(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n574), .B2(new_n575), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n503), .A2(new_n593), .B1(new_n509), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n592), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n512), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n503), .A2(new_n599), .B1(new_n509), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(new_n587), .A2(G54), .ZN(new_n604));
  AND2_X1   g179(.A1(G79), .A2(G543), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n513), .B2(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n606), .B2(new_n512), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n509), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n576), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g190(.A(new_n614), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n580), .B(KEYINPUT75), .Z(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n612), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(new_n549), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n613), .A2(G559), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G323));
  XNOR2_X1  g201(.A(KEYINPUT76), .B(KEYINPUT11), .ZN(new_n627));
  XNOR2_X1  g202(.A(G323), .B(new_n627), .ZN(G282));
  NAND2_X1  g203(.A1(new_n475), .A2(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n475), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n479), .A2(G123), .ZN(new_n636));
  MUX2_X1   g211(.A(G99), .B(G111), .S(G2105), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G2104), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT77), .B(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n633), .A2(new_n634), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT78), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n668), .B2(new_n660), .ZN(new_n669));
  INV_X1    g244(.A(new_n668), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n661), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n661), .A2(new_n664), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n667), .B1(new_n672), .B2(KEYINPUT17), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n632), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT79), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n687), .B(new_n686), .S(new_n679), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT80), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G305), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT84), .B(G1971), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n706), .B2(new_n707), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT83), .B(KEYINPUT34), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  MUX2_X1   g293(.A(G95), .B(G107), .S(G2105), .Z(new_n719));
  AOI22_X1  g294(.A1(new_n479), .A2(G119), .B1(G2104), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G131), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n472), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT81), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G24), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n602), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT82), .B(G1986), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n717), .A2(new_n718), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT36), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n734), .B(new_n736), .Z(new_n737));
  AOI22_X1  g312(.A1(G129), .A2(new_n479), .B1(new_n475), .B2(G141), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G105), .B2(new_n468), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(G29), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT90), .B1(G29), .B2(G32), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n724), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n477), .B2(new_n724), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G171), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT91), .Z(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n753), .B1(new_n757), .B2(G1961), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G162), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n759), .A2(new_n760), .B1(new_n764), .B2(G2090), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G2090), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n704), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n580), .B2(new_n704), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n724), .A2(G33), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n471), .A2(G127), .ZN(new_n773));
  AND2_X1   g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  OAI21_X1  g349(.A(G2105), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n468), .A2(G103), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(new_n475), .B2(G139), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n772), .B1(new_n783), .B2(new_n724), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2072), .ZN(new_n785));
  NOR2_X1   g360(.A1(G27), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G164), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT93), .B(G2078), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(KEYINPUT30), .A2(G28), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT30), .A2(G28), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT31), .B(G11), .Z(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n704), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n704), .B2(G21), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n795), .B1(new_n724), .B2(new_n639), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n800));
  INV_X1    g375(.A(new_n797), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G1966), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n790), .B(new_n803), .C1(new_n804), .C2(new_n756), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n771), .B(new_n805), .C1(new_n760), .C2(new_n759), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n549), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT87), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1341), .ZN(new_n810));
  NOR2_X1   g385(.A1(G4), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n612), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT86), .B(G1348), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G104), .B(G116), .S(G2105), .Z(new_n815));
  AOI22_X1  g390(.A1(new_n479), .A2(G128), .B1(G2104), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G140), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n472), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n724), .A2(G26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT28), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G2067), .Z(new_n823));
  OR2_X1    g398(.A1(new_n812), .A2(new_n813), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n810), .A2(new_n814), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT88), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n737), .A2(new_n766), .A3(new_n806), .A4(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  AOI22_X1  g403(.A1(new_n576), .A2(G93), .B1(new_n587), .B2(G55), .ZN(new_n829));
  OAI21_X1  g404(.A(G67), .B1(new_n506), .B2(new_n505), .ZN(new_n830));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n512), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n543), .A2(new_n544), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G651), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n576), .A2(G81), .B1(new_n587), .B2(G43), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n829), .A4(new_n833), .ZN(new_n840));
  OAI211_X1 g415(.A(G55), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n509), .B2(new_n842), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n545), .A2(new_n548), .B1(new_n843), .B2(new_n832), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n613), .A2(new_n621), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n836), .B1(new_n850), .B2(new_n852), .ZN(G145));
  XOR2_X1   g428(.A(new_n818), .B(KEYINPUT97), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n783), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n490), .A2(new_n497), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n738), .A2(new_n741), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n630), .B(new_n722), .ZN(new_n860));
  MUX2_X1   g435(.A(G106), .B(G118), .S(G2105), .Z(new_n861));
  AOI22_X1  g436(.A1(new_n479), .A2(G130), .B1(G2104), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G142), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n472), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n855), .A2(new_n858), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n859), .A2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n865), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT98), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n871));
  AOI211_X1 g446(.A(new_n871), .B(new_n865), .C1(new_n859), .C2(new_n866), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n477), .B(new_n639), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT96), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n868), .A2(new_n869), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n859), .A2(new_n882), .A3(new_n865), .A4(new_n866), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(new_n879), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g461(.A1(new_n834), .A2(G868), .ZN(new_n887));
  NOR2_X1   g462(.A1(G166), .A2(G305), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n700), .B1(new_n518), .B2(new_n519), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n602), .B(G288), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n888), .B2(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT102), .B1(new_n896), .B2(KEYINPUT42), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  MUX2_X1   g477(.A(KEYINPUT102), .B(new_n897), .S(new_n902), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n612), .A2(new_n568), .A3(new_n579), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT100), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n612), .A2(new_n568), .A3(new_n907), .A4(new_n579), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n612), .B1(new_n568), .B2(new_n579), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g487(.A(KEYINPUT41), .B(new_n910), .C1(new_n906), .C2(new_n908), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n840), .A2(new_n844), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n625), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n906), .B2(new_n908), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n916), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n903), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n887), .B1(new_n920), .B2(G868), .ZN(G295));
  AOI21_X1  g496(.A(new_n887), .B1(new_n920), .B2(G868), .ZN(G331));
  OAI22_X1  g497(.A1(new_n530), .A2(new_n534), .B1(new_n538), .B2(new_n541), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT72), .B(G90), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n576), .A2(new_n924), .B1(new_n587), .B2(G52), .ZN(new_n925));
  NAND3_X1  g500(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n929), .A2(new_n527), .B1(new_n587), .B2(G51), .ZN(new_n930));
  INV_X1    g505(.A(G89), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n574), .B2(new_n575), .ZN(new_n932));
  INV_X1    g507(.A(new_n533), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n513), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n539), .A2(new_n540), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G651), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n925), .A2(new_n930), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n923), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n915), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n840), .A2(new_n923), .A3(new_n937), .A4(new_n844), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n939), .B(new_n940), .Z(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(new_n918), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n923), .A2(new_n937), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n845), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n915), .A2(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(KEYINPUT103), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT104), .B1(new_n914), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n951));
  NOR4_X1   g526(.A1(new_n912), .A2(new_n913), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n901), .B(new_n942), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n879), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n909), .A2(new_n911), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n918), .A2(new_n904), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n949), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n951), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n901), .B1(new_n961), .B2(new_n942), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n914), .A2(new_n941), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n967), .A2(KEYINPUT106), .B1(new_n955), .B2(new_n948), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n914), .A2(new_n969), .A3(new_n941), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n901), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n954), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n965), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n965), .B1(new_n963), .B2(new_n966), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n954), .B2(new_n971), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT107), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n942), .B1(new_n950), .B2(new_n952), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n900), .B2(new_n899), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n966), .A3(new_n879), .A4(new_n953), .ZN(new_n979));
  AND4_X1   g554(.A1(KEYINPUT107), .A2(new_n975), .A3(new_n979), .A4(KEYINPUT44), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n973), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n973), .C1(new_n976), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(G397));
  NAND2_X1  g560(.A1(G303), .A2(G8), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT55), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n500), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT117), .Z(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  NAND2_X1  g568(.A1(G160), .A2(G40), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n495), .B1(new_n487), .B2(new_n489), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT111), .B1(new_n995), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n856), .A2(new_n997), .A3(new_n990), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n992), .A2(new_n993), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1971), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n995), .A2(G1384), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n994), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n500), .A2(new_n990), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n988), .B1(new_n1012), .B2(G8), .ZN(new_n1013));
  AND2_X1   g588(.A1(G160), .A2(G40), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n996), .A3(new_n998), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(G288), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1016), .B(new_n1018), .C1(new_n1017), .C2(G288), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(G1981), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G305), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n592), .B1(KEYINPUT114), .B2(new_n595), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(KEYINPUT114), .B2(new_n595), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(G1981), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1024), .A2(KEYINPUT115), .A3(KEYINPUT49), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n1024), .B2(KEYINPUT49), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1016), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1015), .A2(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(new_n1017), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1019), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1019), .A2(new_n1028), .A3(KEYINPUT118), .A4(new_n1031), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1013), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT50), .B1(new_n996), .B2(new_n998), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1005), .A2(new_n989), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n993), .B(new_n1014), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1011), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1042), .B2(new_n987), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1011), .B2(new_n1040), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT112), .A3(new_n988), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1014), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1053), .A2(new_n1054), .B1(new_n804), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n996), .A2(new_n998), .A3(new_n1007), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n994), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1050), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1048), .A2(G301), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1055), .A2(G2084), .B1(new_n1059), .B2(G1966), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1063), .B2(G286), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1063), .B2(G286), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT125), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1065), .B(new_n1071), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n577), .A2(new_n578), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT57), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1014), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n991), .B(KEYINPUT117), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1049), .A2(new_n1052), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1078), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1015), .A2(G2067), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1055), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n613), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT121), .B(G1996), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1049), .A2(new_n1093), .A3(new_n1052), .A4(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1052), .A2(new_n1008), .A3(new_n1004), .A4(new_n1094), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT122), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1015), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n549), .C1(KEYINPUT123), .C2(KEYINPUT59), .ZN(new_n1102));
  NOR2_X1   g677(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1095), .A2(new_n1097), .B1(new_n1015), .B2(new_n1099), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n623), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1102), .A2(new_n1105), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1083), .A2(new_n1085), .A3(new_n1078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n1090), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1107), .B2(new_n1086), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1087), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1090), .A2(new_n613), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1091), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1092), .B1(new_n1106), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1118), .A2(new_n1054), .A3(G2078), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1004), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G171), .B(KEYINPUT54), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1056), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1061), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1048), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1117), .A2(new_n1124), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1029), .B(KEYINPUT116), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1028), .A2(new_n1017), .A3(new_n710), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1021), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1047), .B2(new_n1032), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  AND4_X1   g705(.A1(KEYINPUT63), .A2(new_n1019), .A3(new_n1028), .A4(new_n1031), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1042), .A2(new_n987), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G286), .A2(new_n1044), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1063), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT119), .B1(new_n1063), .B2(new_n1133), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1131), .B(new_n1132), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1045), .A2(KEYINPUT112), .A3(new_n988), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT112), .B1(new_n1045), .B2(new_n988), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1130), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1047), .A3(KEYINPUT120), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1036), .A2(new_n1047), .A3(new_n1142), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1129), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1075), .A2(new_n1125), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1118), .A2(new_n1014), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n818), .B(G2067), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT109), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(KEYINPUT109), .A3(new_n1152), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n857), .B(G1996), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1153), .B(new_n1154), .C1(new_n1151), .C2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n722), .B(new_n728), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n602), .B(G1986), .Z(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1149), .A2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1150), .A2(G1986), .A3(G290), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n728), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n722), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n818), .A2(G2067), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1150), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OR3_X1    g744(.A1(new_n1150), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT46), .B1(new_n1150), .B2(G1996), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1152), .A2(new_n857), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1170), .A2(new_n1171), .B1(new_n1151), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1164), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1161), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g751(.A1(G401), .A2(new_n459), .ZN(new_n1178));
  AND3_X1   g752(.A1(new_n697), .A2(new_n676), .A3(new_n1178), .ZN(new_n1179));
  NAND4_X1  g753(.A1(new_n885), .A2(new_n972), .A3(new_n964), .A4(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g754(.A(new_n1180), .B(KEYINPUT126), .ZN(G308));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT126), .Z(G225));
endmodule


