//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT68), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n465), .B2(new_n466), .ZN(new_n480));
  AND2_X1   g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n466), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n461), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n485), .A2(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n473), .A2(new_n474), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n461), .A2(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n505), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n502), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n502), .A2(new_n506), .A3(new_n508), .A4(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OR2_X1    g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n518), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  INV_X1    g112(.A(new_n532), .ZN(new_n538));
  NOR2_X1   g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  OAI211_X1 g114(.A(G51), .B(G543), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT7), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n543), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n536), .A2(new_n537), .A3(new_n540), .A4(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(G89), .B1(new_n538), .B2(new_n539), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n540), .A2(new_n545), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT72), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n546), .A2(new_n553), .ZN(G168));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n516), .B2(new_n517), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT73), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n560), .B(new_n557), .C1(new_n549), .C2(new_n555), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(G651), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n516), .A2(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n563));
  INV_X1    g138(.A(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n531), .B2(new_n532), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n563), .A2(G90), .B1(new_n565), .B2(G52), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n562), .A2(new_n566), .ZN(G171));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  INV_X1    g143(.A(G68), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n549), .A2(new_n568), .B1(new_n569), .B2(new_n564), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI221_X1 g147(.A(KEYINPUT74), .B1(new_n569), .B2(new_n564), .C1(new_n549), .C2(new_n568), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G651), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n563), .A2(G81), .B1(new_n565), .B2(G43), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  NAND4_X1  g153(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND4_X1  g156(.A1(G319), .A2(G483), .A3(G661), .A4(new_n581), .ZN(G188));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n549), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n563), .A2(G91), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n565), .A2(G53), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(KEYINPUT9), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT9), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n565), .B2(G53), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n586), .B(new_n587), .C1(new_n589), .C2(new_n591), .ZN(G299));
  NAND2_X1  g167(.A1(new_n562), .A2(new_n566), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n562), .A2(KEYINPUT75), .A3(new_n566), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G301));
  INV_X1    g173(.A(G168), .ZN(G286));
  INV_X1    g174(.A(G166), .ZN(G303));
  INV_X1    g175(.A(G87), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT76), .B1(new_n524), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n563), .A2(new_n603), .A3(G87), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G74), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n516), .A2(new_n606), .A3(new_n517), .ZN(new_n607));
  AOI22_X1  g182(.A1(G49), .A2(new_n565), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(G288));
  INV_X1    g184(.A(G61), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n516), .B2(new_n517), .ZN(new_n611));
  NAND2_X1  g186(.A1(G73), .A2(G543), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT77), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n614), .A2(G73), .A3(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n518), .A2(new_n523), .A3(G86), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n565), .A2(G48), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(G305));
  NAND2_X1  g195(.A1(G72), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G60), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n549), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n515), .B1(new_n623), .B2(KEYINPUT78), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(KEYINPUT78), .B2(new_n623), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n563), .A2(G85), .B1(new_n565), .B2(G47), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(G290));
  XOR2_X1   g202(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G92), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n524), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n563), .A2(G92), .A3(new_n628), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n565), .A2(G54), .ZN(new_n633));
  INV_X1    g208(.A(G66), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n516), .B2(new_n517), .ZN(new_n635));
  AND2_X1   g210(.A1(G79), .A2(G543), .ZN(new_n636));
  OAI21_X1  g211(.A(G651), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n597), .B2(G868), .ZN(G284));
  AOI21_X1  g215(.A(new_n639), .B1(new_n597), .B2(G868), .ZN(G321));
  NOR2_X1   g216(.A1(G299), .A2(G868), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G868), .B2(G168), .ZN(G280));
  XNOR2_X1  g218(.A(G280), .B(KEYINPUT80), .ZN(G297));
  AND4_X1   g219(.A1(new_n633), .A2(new_n631), .A3(new_n637), .A4(new_n632), .ZN(new_n645));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G860), .ZN(G148));
  INV_X1    g222(.A(G868), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n576), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n638), .A2(G559), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(new_n648), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g227(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n653));
  XNOR2_X1  g228(.A(G323), .B(new_n653), .ZN(G282));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n463), .A2(new_n464), .A3(G2105), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT13), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n489), .A2(G135), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n491), .A2(G123), .ZN(new_n661));
  OR2_X1    g236(.A1(G99), .A2(G2105), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n662), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(G2096), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(G2096), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n665), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(G2427), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2430), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT15), .B(G2435), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT14), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2451), .B(G2454), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G14), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G401));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(KEYINPUT85), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(KEYINPUT85), .B2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n685), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n688), .B(new_n690), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n686), .A3(new_n685), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n692), .A2(new_n693), .A3(new_n689), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XNOR2_X1  g275(.A(G2096), .B(G2100), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G227));
  XNOR2_X1  g278(.A(G1971), .B(G1976), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT19), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1956), .B(G2474), .Z(new_n707));
  XOR2_X1   g282(.A(G1961), .B(G1966), .Z(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n714), .B(new_n713), .S(new_n706), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(G1991), .B(G1996), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n717), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n716), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n719), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(G1981), .B(G1986), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n725), .B1(new_n720), .B2(new_n724), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(G229));
  NOR2_X1   g304(.A1(G6), .A2(G16), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT32), .B(G1981), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G23), .ZN(new_n736));
  INV_X1    g311(.A(G288), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n735), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT33), .B(G1976), .Z(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n735), .A2(G22), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G166), .B2(new_n735), .ZN(new_n742));
  INV_X1    g317(.A(G1971), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n744), .C1(new_n738), .C2(new_n739), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT34), .Z(new_n746));
  MUX2_X1   g321(.A(G24), .B(G290), .S(G16), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1986), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n489), .A2(G131), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n491), .A2(G119), .ZN(new_n752));
  OR2_X1    g327(.A1(G95), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT88), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(new_n749), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT35), .B(G1991), .Z(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n748), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n746), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT36), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n735), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n735), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G1966), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT30), .B(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(KEYINPUT31), .A2(G11), .ZN(new_n769));
  NAND2_X1  g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n768), .A2(new_n749), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n664), .B2(new_n749), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n765), .B2(G1966), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  NOR2_X1   g349(.A1(G171), .A2(new_n735), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G5), .B2(new_n735), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n767), .B(new_n773), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n749), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n749), .ZN(new_n780));
  INV_X1    g355(.A(G2090), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n749), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NOR3_X1   g361(.A1(new_n473), .A2(new_n474), .A3(new_n486), .ZN(new_n787));
  AOI21_X1  g362(.A(KEYINPUT69), .B1(new_n465), .B2(new_n466), .ZN(new_n788));
  OAI211_X1 g363(.A(G140), .B(new_n461), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(G128), .B(G2105), .C1(new_n787), .C2(new_n788), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n461), .A2(G116), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT89), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT89), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n789), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n789), .A2(new_n790), .A3(new_n795), .A4(KEYINPUT90), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n786), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G19), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n577), .B2(G16), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1341), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n645), .A2(G16), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G4), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n749), .A2(G33), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(new_n461), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n461), .B1(new_n787), .B2(new_n788), .ZN(new_n819));
  INV_X1    g394(.A(G139), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n815), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n813), .B1(new_n821), .B2(G29), .ZN(new_n822));
  INV_X1    g397(.A(G2072), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n812), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n810), .A2(new_n811), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n735), .A2(G20), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT97), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT23), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G299), .B2(G16), .ZN(new_n831));
  INV_X1    g406(.A(G1956), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G34), .ZN(new_n834));
  AOI21_X1  g409(.A(G29), .B1(new_n834), .B2(KEYINPUT24), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT24), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n483), .B2(new_n749), .ZN(new_n837));
  INV_X1    g412(.A(G2084), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n826), .A2(new_n827), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n831), .A2(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n825), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n784), .A2(new_n805), .A3(new_n808), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n749), .A2(G27), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT94), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G164), .B2(new_n749), .ZN(new_n846));
  INV_X1    g421(.A(G2078), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n489), .A2(G141), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n491), .A2(G129), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT26), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n855), .A2(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n851), .A2(new_n852), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n749), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n749), .B2(G32), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT27), .B(G1996), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n774), .B2(new_n776), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR4_X1   g445(.A1(new_n843), .A2(new_n849), .A3(new_n850), .A4(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n763), .A2(new_n778), .A3(new_n871), .ZN(G311));
  NAND3_X1  g447(.A1(new_n763), .A2(new_n778), .A3(new_n871), .ZN(G150));
  NAND2_X1  g448(.A1(new_n645), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT38), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n515), .ZN(new_n877));
  INV_X1    g452(.A(G93), .ZN(new_n878));
  INV_X1    g453(.A(G55), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n524), .A2(new_n878), .B1(new_n526), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n576), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n875), .B(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  INV_X1    g459(.A(G860), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n881), .A2(new_n885), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(G145));
  XNOR2_X1  g465(.A(new_n657), .B(KEYINPUT102), .ZN(new_n891));
  INV_X1    g466(.A(G142), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n819), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n489), .A2(new_n894), .A3(G142), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(G118), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(G2105), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n491), .B2(G130), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n756), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n756), .B1(new_n896), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n891), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n896), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n757), .ZN(new_n906));
  INV_X1    g481(.A(new_n891), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n509), .B1(new_n798), .B2(new_n800), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n798), .A2(new_n509), .A3(new_n800), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n863), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n798), .A2(new_n509), .A3(new_n800), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n862), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  INV_X1    g490(.A(new_n821), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT99), .B1(new_n916), .B2(KEYINPUT100), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n916), .A2(KEYINPUT99), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n913), .A2(new_n915), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(KEYINPUT103), .B(new_n909), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n664), .B(KEYINPUT98), .Z(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G160), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n664), .B(KEYINPUT98), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n483), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n495), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n925), .A3(G162), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n913), .A2(new_n915), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n917), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n902), .A2(new_n903), .A3(new_n891), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n907), .B1(new_n906), .B2(new_n901), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT103), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n904), .A2(new_n936), .A3(new_n908), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n921), .A2(new_n929), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n929), .B1(new_n921), .B2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g522(.A1(new_n877), .A2(new_n880), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n648), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n882), .B(new_n650), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT104), .B1(new_n645), .B2(G299), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n645), .A2(G299), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n588), .B(KEYINPUT9), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n586), .A2(new_n587), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n638), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n954), .A3(new_n638), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n645), .B2(G299), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n957), .A2(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n952), .A2(new_n959), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n950), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G166), .A2(G290), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n625), .B(new_n626), .C1(new_n522), .C2(new_n528), .ZN(new_n967));
  NAND2_X1  g542(.A1(G288), .A2(new_n731), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n737), .A2(G305), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n966), .A2(new_n967), .B1(new_n969), .B2(new_n968), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n965), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n949), .B1(new_n974), .B2(new_n648), .ZN(G295));
  OAI21_X1  g550(.A(new_n949), .B1(new_n974), .B2(new_n648), .ZN(G331));
  INV_X1    g551(.A(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n957), .A2(new_n958), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n960), .A2(new_n959), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n576), .B(new_n948), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n595), .A2(G168), .A3(new_n596), .ZN(new_n982));
  NAND4_X1  g557(.A1(G171), .A2(KEYINPUT106), .A3(new_n546), .A4(new_n553), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G168), .B2(new_n593), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n882), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n980), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n986), .A2(new_n963), .A3(new_n988), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n977), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n991), .B2(KEYINPUT107), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n987), .A2(new_n882), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n987), .A2(new_n882), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n961), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n986), .A2(new_n963), .A3(new_n988), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n972), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n958), .B1(new_n986), .B2(new_n988), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n977), .B1(new_n957), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n964), .B2(new_n1001), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n992), .A2(new_n999), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n941), .B1(new_n997), .B2(new_n998), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n989), .A2(new_n990), .A3(new_n977), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT107), .B(new_n972), .C1(new_n995), .C2(new_n996), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(new_n1000), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n992), .A2(new_n999), .A3(new_n1003), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1008), .A2(new_n1000), .B1(new_n1010), .B2(KEYINPUT43), .ZN(new_n1011));
  MUX2_X1   g586(.A(new_n1009), .B(new_n1011), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g587(.A(new_n802), .B(G2067), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n862), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n756), .B(new_n759), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(G290), .B(G1986), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n475), .A2(new_n476), .A3(new_n468), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n476), .B1(new_n475), .B2(new_n468), .ZN(new_n1023));
  OAI211_X1 g598(.A(G40), .B(new_n482), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT108), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n478), .A2(new_n1026), .A3(G40), .A4(new_n482), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n509), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1021), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1030), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1025), .A2(new_n1038), .A3(new_n1027), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n499), .A2(new_n501), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n497), .B1(new_n473), .B2(new_n474), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT4), .B1(new_n485), .B2(new_n507), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT70), .B1(new_n1046), .B2(new_n508), .ZN(new_n1047));
  INV_X1    g622(.A(new_n512), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1041), .B(new_n1029), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1956), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n513), .B2(new_n1029), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1025), .A2(new_n1027), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1035), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n513), .A2(new_n1029), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1031), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1025), .A2(new_n1027), .A3(new_n1052), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1054), .ZN(new_n1061));
  AOI211_X1 g636(.A(KEYINPUT50), .B(G1384), .C1(new_n511), .C2(new_n512), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n832), .B1(new_n1039), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(KEYINPUT119), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n953), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(G299), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1057), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(KEYINPUT50), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n509), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1025), .A2(new_n1027), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1041), .B1(new_n513), .B2(new_n1029), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1025), .A2(new_n1027), .A3(new_n1071), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT118), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n811), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1030), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1025), .A2(new_n1079), .A3(new_n1027), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(G2067), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1061), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n645), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1069), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1061), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1084), .B2(KEYINPUT121), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1069), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1067), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT120), .B(G1996), .Z(new_n1095));
  NOR3_X1   g670(.A1(new_n1051), .A2(new_n1053), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1080), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n577), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT59), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1102), .B(new_n577), .C1(new_n1096), .C2(new_n1099), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1092), .A2(new_n1094), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n638), .A2(KEYINPUT122), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n638), .A2(KEYINPUT122), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1083), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1082), .A2(new_n1107), .A3(new_n1106), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1082), .A2(new_n1107), .B1(KEYINPUT122), .B2(new_n638), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1086), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n1115));
  INV_X1    g690(.A(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(G166), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT55), .B(G8), .C1(new_n522), .C2(new_n528), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n743), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1049), .A2(new_n1025), .A3(new_n1027), .A4(new_n1038), .ZN(new_n1122));
  AOI21_X1  g697(.A(G2090), .B1(new_n1122), .B2(KEYINPUT115), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1039), .A2(new_n1062), .A3(KEYINPUT115), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1119), .B1(new_n1125), .B2(new_n1116), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n603), .B1(new_n563), .B2(G87), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n603), .A2(new_n518), .A3(new_n523), .A4(G87), .ZN(new_n1128));
  OAI211_X1 g703(.A(G1976), .B(new_n608), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT113), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n605), .A2(new_n1131), .A3(G1976), .A4(new_n608), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(new_n1080), .A3(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT52), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1133), .A2(new_n1080), .A3(G8), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(G305), .A2(G1981), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1981), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n617), .A2(new_n1141), .A3(new_n618), .A4(new_n619), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT49), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1139), .A3(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n1151), .A3(G8), .A4(new_n1080), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1135), .A2(new_n1138), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT116), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT116), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1135), .A2(new_n1152), .A3(new_n1155), .A4(new_n1138), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT112), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1117), .A2(new_n1158), .A3(new_n1118), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT111), .B1(new_n1162), .B2(new_n781), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1070), .A2(new_n1072), .A3(KEYINPUT111), .A4(new_n781), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1120), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1161), .B(G8), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1126), .A2(new_n1157), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT51), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n838), .ZN(new_n1170));
  INV_X1    g745(.A(G1966), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1025), .A2(new_n1032), .A3(new_n1027), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1170), .A2(new_n1175), .A3(G168), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT51), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1116), .B1(KEYINPUT123), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1169), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(G8), .A3(G286), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1176), .A2(new_n1178), .A3(new_n1169), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1051), .A2(new_n1053), .A3(G2078), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT53), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1074), .A2(new_n774), .A3(new_n1077), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1174), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1172), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1187), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1188), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1193));
  OAI211_X1 g768(.A(G301), .B(new_n1186), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1024), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1196), .A2(new_n1052), .A3(new_n1190), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1185), .B2(KEYINPUT53), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1187), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1074), .A2(new_n1077), .A3(KEYINPUT125), .A4(new_n774), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(KEYINPUT54), .B1(new_n1202), .B2(new_n593), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1167), .B(new_n1184), .C1(new_n1195), .C2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n597), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1202), .A2(G301), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT54), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1114), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1206), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1183), .A2(new_n1182), .ZN(new_n1211));
  OAI21_X1  g786(.A(KEYINPUT62), .B1(new_n1211), .B2(new_n1179), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1180), .A2(new_n1213), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1210), .A2(new_n1212), .A3(new_n1214), .A4(new_n1167), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n1116), .B(G286), .C1(new_n1170), .C2(new_n1175), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1126), .A2(new_n1157), .A3(new_n1166), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(G8), .B1(new_n1165), .B2(new_n1163), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n1119), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1153), .A2(new_n1218), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1221), .A2(new_n1166), .A3(new_n1216), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1166), .A2(new_n1153), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1152), .A2(new_n1136), .A3(new_n737), .ZN(new_n1226));
  AOI211_X1 g801(.A(new_n1116), .B(new_n1097), .C1(new_n1226), .C2(new_n1142), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1215), .A2(new_n1224), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1034), .B1(new_n1209), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1033), .A2(new_n1014), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1231), .B(KEYINPUT46), .Z(new_n1232));
  INV_X1    g807(.A(new_n1033), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1013), .B2(new_n863), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT47), .Z(new_n1236));
  NOR3_X1   g811(.A1(new_n1233), .A2(G1986), .A3(G290), .ZN(new_n1237));
  XOR2_X1   g812(.A(new_n1237), .B(KEYINPUT48), .Z(new_n1238));
  OAI21_X1  g813(.A(new_n1238), .B1(new_n1233), .B2(new_n1019), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n757), .A2(new_n759), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1240), .B(KEYINPUT126), .ZN(new_n1241));
  OAI22_X1  g816(.A1(new_n1016), .A2(new_n1241), .B1(G2067), .B2(new_n803), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1242), .A2(new_n1033), .ZN(new_n1243));
  AND3_X1   g818(.A1(new_n1236), .A2(new_n1239), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1230), .A2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1247));
  OAI211_X1 g821(.A(new_n702), .B(G319), .C1(new_n683), .C2(new_n682), .ZN(new_n1248));
  NAND2_X1  g822(.A1(new_n720), .A2(new_n724), .ZN(new_n1249));
  INV_X1    g823(.A(new_n725), .ZN(new_n1250));
  NAND2_X1  g824(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1248), .B1(new_n1251), .B2(new_n726), .ZN(new_n1252));
  OAI21_X1  g826(.A(new_n1252), .B1(new_n942), .B2(new_n944), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n991), .A2(KEYINPUT107), .ZN(new_n1254));
  INV_X1    g828(.A(new_n1006), .ZN(new_n1255));
  NAND4_X1  g829(.A1(new_n1254), .A2(new_n1255), .A3(new_n941), .A4(new_n999), .ZN(new_n1256));
  INV_X1    g830(.A(new_n1000), .ZN(new_n1257));
  NAND2_X1  g831(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g832(.A(new_n1247), .B(new_n1253), .C1(new_n1258), .C2(new_n1004), .ZN(new_n1259));
  INV_X1    g833(.A(new_n1253), .ZN(new_n1260));
  AOI21_X1  g834(.A(KEYINPUT127), .B1(new_n1009), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g835(.A1(new_n1259), .A2(new_n1261), .ZN(G308));
  NAND2_X1  g836(.A1(new_n1009), .A2(new_n1260), .ZN(new_n1263));
  NAND2_X1  g837(.A1(new_n1263), .A2(new_n1247), .ZN(new_n1264));
  NAND3_X1  g838(.A1(new_n1009), .A2(new_n1260), .A3(KEYINPUT127), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n1264), .A2(new_n1265), .ZN(G225));
endmodule


