

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X2 U320 ( .A(n440), .B(KEYINPUT48), .ZN(n546) );
  XNOR2_X1 U321 ( .A(n427), .B(n426), .ZN(n573) );
  XNOR2_X1 U322 ( .A(n421), .B(n420), .ZN(n425) );
  XNOR2_X1 U323 ( .A(n442), .B(KEYINPUT54), .ZN(n443) );
  XNOR2_X1 U324 ( .A(n395), .B(n288), .ZN(n396) );
  XOR2_X1 U325 ( .A(n394), .B(n393), .Z(n288) );
  XOR2_X1 U326 ( .A(KEYINPUT45), .B(n404), .Z(n289) );
  XNOR2_X1 U327 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U328 ( .A(n410), .B(n409), .ZN(n413) );
  INV_X1 U329 ( .A(n416), .ZN(n419) );
  INV_X1 U330 ( .A(KEYINPUT119), .ZN(n442) );
  XNOR2_X1 U331 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U332 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U333 ( .A(KEYINPUT36), .ZN(n402) );
  XNOR2_X1 U334 ( .A(n402), .B(KEYINPUT96), .ZN(n403) );
  XNOR2_X1 U335 ( .A(n432), .B(n403), .ZN(n582) );
  NOR2_X2 U336 ( .A1(n460), .A2(n448), .ZN(n560) );
  XNOR2_X1 U337 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n423) );
  XOR2_X1 U340 ( .A(G127GAT), .B(KEYINPUT0), .Z(n291) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(G134GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n332) );
  XOR2_X1 U343 ( .A(n423), .B(n332), .Z(n293) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U346 ( .A(n294), .B(G176GAT), .Z(n298) );
  XOR2_X1 U347 ( .A(G183GAT), .B(KEYINPUT18), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n341) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(n341), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n306) );
  XOR2_X1 U352 ( .A(G190GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G43GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(n304), .B(n303), .Z(n305) );
  XOR2_X2 U359 ( .A(n306), .B(n305), .Z(n530) );
  INV_X1 U360 ( .A(n530), .ZN(n460) );
  XNOR2_X1 U361 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n307), .B(KEYINPUT2), .ZN(n331) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n392) );
  XOR2_X1 U364 ( .A(n331), .B(n392), .Z(n309) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U367 ( .A(n310), .B(KEYINPUT23), .Z(n312) );
  XOR2_X1 U368 ( .A(G141GAT), .B(G22GAT), .Z(n351) );
  XNOR2_X1 U369 ( .A(n351), .B(KEYINPUT24), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U371 ( .A(G204GAT), .B(KEYINPUT85), .Z(n314) );
  XNOR2_X1 U372 ( .A(KEYINPUT22), .B(KEYINPUT84), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U374 ( .A(n316), .B(n315), .Z(n322) );
  XOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n349) );
  XOR2_X1 U378 ( .A(G78GAT), .B(G148GAT), .Z(n320) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n410) );
  XNOR2_X1 U381 ( .A(n349), .B(n410), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n469) );
  XOR2_X1 U383 ( .A(KEYINPUT1), .B(KEYINPUT86), .Z(n324) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(G57GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n340) );
  XOR2_X1 U386 ( .A(G148GAT), .B(G120GAT), .Z(n326) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(G141GAT), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U389 ( .A(G162GAT), .B(G85GAT), .Z(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n336) );
  XNOR2_X1 U391 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n329), .B(KEYINPUT87), .ZN(n330) );
  XOR2_X1 U393 ( .A(n330), .B(KEYINPUT5), .Z(n334) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n338) );
  NAND2_X1 U397 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n518) );
  XOR2_X1 U400 ( .A(G169GAT), .B(G8GAT), .Z(n352) );
  XNOR2_X1 U401 ( .A(n352), .B(n341), .ZN(n347) );
  XOR2_X1 U402 ( .A(G36GAT), .B(G190GAT), .Z(n386) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G92GAT), .Z(n343) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n416) );
  XOR2_X1 U406 ( .A(n386), .B(n416), .Z(n345) );
  NAND2_X1 U407 ( .A1(G226GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n520) );
  XNOR2_X1 U411 ( .A(KEYINPUT118), .B(n520), .ZN(n441) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G1GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n350), .B(KEYINPUT70), .ZN(n373) );
  XNOR2_X1 U414 ( .A(n351), .B(n373), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n359) );
  XOR2_X1 U416 ( .A(G29GAT), .B(G43GAT), .Z(n355) );
  XNOR2_X1 U417 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n399) );
  XOR2_X1 U419 ( .A(n399), .B(KEYINPUT69), .Z(n357) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U422 ( .A(n359), .B(n358), .Z(n367) );
  XOR2_X1 U423 ( .A(G197GAT), .B(G113GAT), .Z(n361) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(G36GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U426 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n363) );
  XNOR2_X1 U427 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n367), .B(n366), .Z(n505) );
  INV_X1 U431 ( .A(n505), .ZN(n570) );
  XOR2_X1 U432 ( .A(G211GAT), .B(G127GAT), .Z(n369) );
  XNOR2_X1 U433 ( .A(G183GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U435 ( .A(KEYINPUT13), .B(G57GAT), .Z(n417) );
  XOR2_X1 U436 ( .A(n370), .B(n417), .Z(n372) );
  XNOR2_X1 U437 ( .A(G22GAT), .B(G78GAT), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U439 ( .A(n373), .B(KEYINPUT12), .Z(n375) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U442 ( .A(n377), .B(n376), .Z(n385) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n379) );
  XNOR2_X1 U444 ( .A(G155GAT), .B(KEYINPUT80), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U446 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n381) );
  XNOR2_X1 U447 ( .A(G8GAT), .B(G64GAT), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U450 ( .A(n385), .B(n384), .Z(n577) );
  INV_X1 U451 ( .A(n577), .ZN(n489) );
  XOR2_X1 U452 ( .A(G99GAT), .B(G85GAT), .Z(n422) );
  XOR2_X1 U453 ( .A(n422), .B(n386), .Z(n388) );
  NAND2_X1 U454 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n397) );
  XOR2_X1 U456 ( .A(G92GAT), .B(G106GAT), .Z(n390) );
  XNOR2_X1 U457 ( .A(G134GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n395) );
  XOR2_X1 U460 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n394) );
  XNOR2_X1 U461 ( .A(KEYINPUT76), .B(KEYINPUT9), .ZN(n393) );
  XOR2_X1 U462 ( .A(n398), .B(KEYINPUT11), .Z(n401) );
  XNOR2_X1 U463 ( .A(n399), .B(KEYINPUT10), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n432) );
  NOR2_X1 U465 ( .A1(n489), .A2(n582), .ZN(n404) );
  NOR2_X1 U466 ( .A1(n570), .A2(n289), .ZN(n428) );
  XOR2_X1 U467 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n406) );
  XNOR2_X1 U468 ( .A(KEYINPUT31), .B(KEYINPUT72), .ZN(n405) );
  XOR2_X1 U469 ( .A(n406), .B(n405), .Z(n427) );
  NAND2_X1 U470 ( .A1(G230GAT), .A2(G233GAT), .ZN(n408) );
  INV_X1 U471 ( .A(KEYINPUT32), .ZN(n407) );
  INV_X1 U472 ( .A(n413), .ZN(n411) );
  NAND2_X1 U473 ( .A1(n411), .A2(KEYINPUT75), .ZN(n415) );
  INV_X1 U474 ( .A(KEYINPUT75), .ZN(n412) );
  NAND2_X1 U475 ( .A1(n413), .A2(n412), .ZN(n414) );
  NAND2_X1 U476 ( .A1(n415), .A2(n414), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n417), .B(KEYINPUT71), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U480 ( .A1(n428), .A2(n573), .ZN(n439) );
  XOR2_X1 U481 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n429) );
  XOR2_X1 U482 ( .A(n573), .B(n429), .Z(n559) );
  AND2_X1 U483 ( .A1(n570), .A2(n559), .ZN(n431) );
  XNOR2_X1 U484 ( .A(KEYINPUT107), .B(KEYINPUT46), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n434) );
  NOR2_X1 U486 ( .A1(n432), .A2(n577), .ZN(n433) );
  AND2_X1 U487 ( .A1(n434), .A2(n433), .ZN(n437) );
  XOR2_X1 U488 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n435) );
  XNOR2_X1 U489 ( .A(KEYINPUT47), .B(n435), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U491 ( .A1(n439), .A2(n438), .ZN(n440) );
  NAND2_X1 U492 ( .A1(n441), .A2(n546), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U494 ( .A1(n518), .A2(n445), .ZN(n446) );
  XNOR2_X1 U495 ( .A(n446), .B(KEYINPUT65), .ZN(n568) );
  NOR2_X1 U496 ( .A1(n469), .A2(n568), .ZN(n447) );
  XNOR2_X1 U497 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NAND2_X1 U498 ( .A1(n560), .A2(n432), .ZN(n451) );
  XOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n449) );
  NAND2_X1 U500 ( .A1(n560), .A2(n570), .ZN(n453) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n453), .B(n452), .ZN(G1348GAT) );
  NAND2_X1 U503 ( .A1(n577), .A2(n560), .ZN(n455) );
  XNOR2_X1 U504 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  NAND2_X1 U506 ( .A1(n570), .A2(n573), .ZN(n491) );
  NOR2_X1 U507 ( .A1(n432), .A2(n489), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n456), .B(KEYINPUT16), .ZN(n476) );
  AND2_X1 U509 ( .A1(n520), .A2(n530), .ZN(n457) );
  NOR2_X1 U510 ( .A1(n469), .A2(n457), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT91), .ZN(n466) );
  XOR2_X1 U513 ( .A(KEYINPUT26), .B(KEYINPUT89), .Z(n462) );
  NAND2_X1 U514 ( .A1(n469), .A2(n460), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n569) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(n520), .ZN(n470) );
  INV_X1 U517 ( .A(n470), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n569), .A2(n463), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT90), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT92), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n518), .A2(n468), .ZN(n474) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT28), .ZN(n525) );
  INV_X1 U524 ( .A(n525), .ZN(n472) );
  NAND2_X1 U525 ( .A1(n518), .A2(n470), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT88), .B(n471), .Z(n545) );
  NAND2_X1 U527 ( .A1(n472), .A2(n545), .ZN(n532) );
  NOR2_X1 U528 ( .A1(n530), .A2(n532), .ZN(n473) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n487) );
  INV_X1 U530 ( .A(n487), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n507) );
  NOR2_X1 U532 ( .A1(n491), .A2(n507), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n518), .A2(n484), .ZN(n479) );
  XOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT34), .Z(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT93), .B(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n520), .A2(n484), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U540 ( .A1(n484), .A2(n530), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n483), .ZN(G1326GAT) );
  XOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT95), .Z(n486) );
  NAND2_X1 U544 ( .A1(n484), .A2(n525), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U547 ( .A1(n487), .A2(n582), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n490), .Z(n516) );
  NOR2_X1 U550 ( .A1(n491), .A2(n516), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT38), .ZN(n499) );
  NAND2_X1 U552 ( .A1(n499), .A2(n518), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT97), .Z(n496) );
  NAND2_X1 U555 ( .A1(n499), .A2(n520), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n530), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n501) );
  NAND2_X1 U561 ( .A1(n499), .A2(n525), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT102), .ZN(n504) );
  XOR2_X1 U566 ( .A(KEYINPUT101), .B(n504), .Z(n509) );
  NAND2_X1 U567 ( .A1(n505), .A2(n559), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(KEYINPUT100), .ZN(n517) );
  NOR2_X1 U569 ( .A1(n517), .A2(n507), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n518), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n520), .A2(n512), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n512), .A2(n530), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U577 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NOR2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(KEYINPUT104), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT105), .Z(n524) );
  NAND2_X1 U587 ( .A1(n526), .A2(n530), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n528) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n546), .ZN(n531) );
  NOR2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n540), .A2(n570), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n535) );
  NAND2_X1 U598 ( .A1(n540), .A2(n559), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT110), .Z(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n577), .A2(n540), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n432), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT113), .Z(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT115), .Z(n550) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n547), .A2(n569), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT114), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n570), .A2(n556), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n559), .A2(n556), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n556), .A2(n577), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  XOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT117), .Z(n558) );
  NAND2_X1 U624 ( .A1(n432), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT121), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(n567), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n578), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U639 ( .A(n578), .ZN(n581) );
  OR2_X1 U640 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

