//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT0), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n192), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(KEYINPUT64), .B2(new_n194), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n190), .A2(new_n195), .B1(new_n193), .B2(new_n187), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n187), .A2(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n187), .A2(new_n200), .A3(G128), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  OR3_X1    g016(.A1(new_n200), .A2(new_n202), .A3(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(G125), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G224), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(new_n206), .B2(G953), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n205), .B(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G113), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G116), .B(G119), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT5), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n214), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G104), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G107), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n225), .A3(G104), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n234), .A3(new_n228), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n223), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n239), .B(KEYINPUT8), .Z(new_n240));
  INV_X1    g054(.A(new_n237), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n213), .B1(new_n219), .B2(new_n217), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n221), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n208), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n241), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n224), .B1(new_n235), .B2(KEYINPUT82), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(KEYINPUT82), .B2(new_n235), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT4), .A3(new_n236), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n216), .A2(new_n220), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n221), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n251), .C1(KEYINPUT4), .C2(new_n248), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n252), .A3(new_n239), .ZN(new_n253));
  AOI21_X1  g067(.A(G902), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n246), .A2(new_n252), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n239), .B(KEYINPUT85), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n257), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n253), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n257), .A2(KEYINPUT6), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n206), .A2(G953), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT87), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n205), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n254), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G210), .B1(G237), .B2(G902), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(new_n254), .C1(new_n263), .C2(new_n267), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G214), .B1(G237), .B2(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G113), .B(G122), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(new_n227), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT16), .ZN(new_n279));
  INV_X1    g093(.A(G140), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G125), .ZN(new_n281));
  XNOR2_X1  g095(.A(G125), .B(G140), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n284), .A2(new_n202), .ZN(new_n285));
  NOR2_X1   g099(.A1(G237), .A2(G953), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n286), .A2(G143), .A3(G214), .ZN(new_n287));
  AOI21_X1  g101(.A(G143), .B1(new_n286), .B2(G214), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G131), .B1(new_n287), .B2(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n282), .B(KEYINPUT19), .Z(new_n294));
  OAI211_X1 g108(.A(new_n285), .B(new_n293), .C1(G146), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n202), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n283), .A2(G146), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT18), .A2(G131), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n296), .A2(new_n297), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n289), .B2(new_n298), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n278), .B1(new_n301), .B2(KEYINPUT88), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(KEYINPUT88), .B2(new_n301), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n284), .B(G146), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT17), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(new_n292), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n293), .A2(KEYINPUT17), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n278), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G475), .A2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT20), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(KEYINPUT89), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n308), .B2(new_n315), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G475), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G122), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G107), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n210), .A2(KEYINPUT14), .A3(G122), .ZN(new_n323));
  OAI211_X1 g137(.A(G107), .B(new_n323), .C1(new_n321), .C2(KEYINPUT14), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT92), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n192), .A2(G143), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n192), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(KEYINPUT65), .A2(G134), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n334), .ZN(new_n336));
  AOI211_X1 g150(.A(new_n322), .B(new_n325), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n320), .A2(new_n225), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n322), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n328), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n327), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n342), .A2(KEYINPUT91), .B1(new_n326), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(KEYINPUT91), .B2(new_n342), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n339), .B1(new_n344), .B2(G134), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT9), .B(G234), .ZN(new_n346));
  INV_X1    g160(.A(G217), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n346), .A2(new_n347), .A3(G953), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OR3_X1    g163(.A1(new_n337), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n337), .B2(new_n345), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G902), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G478), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(KEYINPUT15), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT93), .A2(G952), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT93), .A2(G952), .ZN(new_n360));
  AOI21_X1  g174(.A(G953), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G234), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G953), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n353), .B(new_n365), .C1(G234), .C2(G237), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT21), .B(G898), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n319), .A2(new_n357), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G469), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT12), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n237), .B(new_n204), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT11), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(new_n331), .A3(G137), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n332), .A2(G137), .A3(new_n333), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n290), .ZN(new_n377));
  AOI21_X1  g191(.A(G137), .B1(new_n332), .B2(new_n333), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT66), .B1(new_n378), .B2(KEYINPUT11), .ZN(new_n379));
  INV_X1    g193(.A(G137), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT65), .A2(G134), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT65), .A2(G134), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT66), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n374), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n375), .B(new_n377), .C1(new_n379), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n375), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n383), .A2(new_n384), .A3(new_n374), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n384), .B1(new_n383), .B2(new_n374), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n376), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(G131), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n372), .B1(new_n373), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  INV_X1    g207(.A(new_n204), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n237), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(G131), .ZN(new_n396));
  INV_X1    g210(.A(new_n377), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n387), .B(new_n397), .C1(new_n388), .C2(new_n389), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(KEYINPUT12), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n392), .A2(new_n393), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n393), .B1(new_n392), .B2(new_n400), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n365), .A2(G227), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n241), .A2(new_n204), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n249), .B(new_n196), .C1(KEYINPUT4), .C2(new_n248), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n204), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n406), .B1(new_n412), .B2(new_n399), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n401), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n412), .A2(new_n399), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n399), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n371), .B(new_n353), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n392), .A2(new_n400), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(new_n399), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n406), .A3(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(G469), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n371), .A2(new_n353), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G221), .B1(new_n346), .B2(G902), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT80), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT81), .Z(new_n429));
  AND2_X1   g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n276), .A2(new_n370), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G217), .B1(new_n362), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n192), .A2(G119), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n212), .A2(G128), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT24), .B(G110), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n434), .A2(new_n437), .ZN(new_n442));
  OAI22_X1  g256(.A1(new_n439), .A2(G110), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n285), .A2(new_n443), .A3(new_n296), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(G110), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n304), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n365), .A2(G221), .A3(G234), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT22), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(G137), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n448), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n353), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT25), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT77), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n433), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n454), .A2(KEYINPUT77), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n457), .A2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n362), .B2(G217), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(G472), .A2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n399), .A2(new_n196), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n380), .A2(G134), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n378), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n383), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT67), .A3(G131), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n398), .A3(new_n204), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(KEYINPUT30), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n398), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n394), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n398), .A3(KEYINPUT68), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n479), .A2(new_n480), .B1(new_n399), .B2(new_n196), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n251), .B(new_n476), .C1(new_n481), .C2(KEYINPUT30), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n251), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n466), .A3(new_n475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n286), .A2(G210), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT27), .Z(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT26), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n224), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT71), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n482), .A2(new_n492), .A3(new_n485), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT31), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT31), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n251), .B(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n475), .B1(new_n391), .B2(new_n197), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT73), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n466), .A2(new_n502), .A3(new_n475), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT28), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g319(.A(new_n251), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n481), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT67), .B1(new_n472), .B2(G131), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n469), .B(new_n290), .C1(new_n383), .C2(new_n471), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n478), .B1(new_n386), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n204), .A3(new_n480), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n466), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT72), .A3(new_n251), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n485), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n504), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT74), .B1(new_n516), .B2(new_n489), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n506), .B1(new_n512), .B2(new_n466), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n485), .B1(new_n518), .B2(KEYINPUT72), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n481), .A2(new_n505), .A3(new_n506), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n504), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n524));
  INV_X1    g338(.A(new_n489), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n498), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n498), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n465), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n516), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n504), .A2(KEYINPUT76), .ZN(new_n537));
  INV_X1    g351(.A(new_n485), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n484), .B1(new_n466), .B2(new_n475), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(KEYINPUT76), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n489), .B(new_n536), .C1(new_n542), .C2(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n482), .A2(new_n485), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(new_n489), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n545), .B2(new_n535), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n534), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n548));
  AOI211_X1 g362(.A(KEYINPUT74), .B(new_n489), .C1(new_n521), .C2(new_n522), .ZN(new_n549));
  INV_X1    g363(.A(new_n497), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT75), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n498), .A2(new_n527), .A3(new_n528), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n465), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n532), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n547), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI211_X1 g372(.A(KEYINPUT79), .B(new_n464), .C1(new_n533), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT79), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n529), .B2(new_n530), .ZN(new_n561));
  INV_X1    g375(.A(new_n547), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(KEYINPUT32), .ZN(new_n564));
  INV_X1    g378(.A(new_n464), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n432), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  OAI21_X1  g382(.A(new_n353), .B1(new_n529), .B2(new_n530), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G472), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n531), .A3(new_n430), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n464), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n319), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n355), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n351), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n352), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n352), .A2(new_n579), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(G478), .B1(new_n352), .B2(new_n353), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n369), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n276), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n573), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n313), .B2(KEYINPUT20), .ZN(new_n593));
  INV_X1    g407(.A(new_n313), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT20), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(KEYINPUT95), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n593), .B(new_n596), .C1(new_n595), .C2(new_n594), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n318), .A3(new_n357), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n588), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n572), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G107), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  INV_X1    g416(.A(new_n571), .ZN(new_n603));
  INV_X1    g417(.A(new_n451), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n448), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n460), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n459), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n370), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n275), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  NAND2_X1  g427(.A1(new_n430), .A2(new_n608), .ZN(new_n614));
  INV_X1    g428(.A(new_n364), .ZN(new_n615));
  INV_X1    g429(.A(G900), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n366), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n317), .B2(G475), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n597), .A2(new_n357), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n564), .A2(new_n276), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n564), .A2(new_n623), .A3(new_n276), .A4(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XOR2_X1   g440(.A(new_n617), .B(KEYINPUT39), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n430), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT40), .Z(new_n629));
  XOR2_X1   g443(.A(new_n273), .B(KEYINPUT38), .Z(new_n630));
  NAND3_X1  g444(.A1(new_n319), .A2(new_n357), .A3(new_n274), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n608), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n494), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n525), .B1(new_n538), .B2(new_n539), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n534), .B1(new_n635), .B2(new_n353), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n555), .B2(new_n557), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n533), .A2(new_n637), .A3(KEYINPUT97), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT97), .B1(new_n533), .B2(new_n637), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n629), .B(new_n632), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G143), .ZN(G45));
  INV_X1    g455(.A(new_n614), .ZN(new_n642));
  INV_X1    g456(.A(new_n617), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n319), .B(new_n643), .C1(new_n582), .C2(new_n583), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n564), .A2(new_n276), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  OR2_X1    g461(.A1(new_n414), .A2(new_n417), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n353), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G469), .ZN(new_n650));
  INV_X1    g464(.A(new_n428), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n418), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n588), .A2(new_n586), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n564), .A3(new_n565), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G113), .ZN(G15));
  INV_X1    g470(.A(new_n652), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n564), .A2(new_n599), .A3(new_n565), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G116), .ZN(G18));
  NOR3_X1   g473(.A1(new_n609), .A2(new_n275), .A3(new_n652), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n564), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G119), .ZN(G21));
  INV_X1    g476(.A(new_n273), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n652), .A2(new_n663), .A3(new_n631), .A4(new_n369), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n498), .B1(new_n489), .B2(new_n542), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n465), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n570), .A2(new_n664), .A3(new_n565), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G122), .ZN(G24));
  NOR3_X1   g483(.A1(new_n652), .A2(new_n275), .A3(new_n644), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n570), .A2(new_n608), .A3(new_n666), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G125), .ZN(G27));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n423), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT99), .A4(G469), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n418), .A2(new_n674), .A3(new_n425), .A4(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n677), .A3(new_n651), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n677), .B1(new_n676), .B2(new_n651), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n271), .A2(new_n274), .A3(new_n272), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n678), .A2(new_n644), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n683), .B(new_n464), .C1(new_n533), .C2(new_n558), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT102), .B1(new_n564), .B2(new_n565), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n564), .A2(new_n565), .A3(new_n681), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n290), .ZN(G33));
  AOI21_X1  g508(.A(new_n464), .B1(new_n533), .B2(new_n558), .ZN(new_n695));
  INV_X1    g509(.A(new_n619), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G134), .ZN(G36));
  NOR2_X1   g513(.A1(new_n584), .A2(new_n319), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT43), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n608), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n570), .A2(new_n531), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT106), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n421), .A2(new_n422), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(G469), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n709), .A2(KEYINPUT104), .A3(G469), .A4(new_n710), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n424), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n418), .B1(new_n715), .B2(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n651), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n627), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n704), .B2(new_n705), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n702), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n703), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n680), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n707), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT107), .B(G137), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G39));
  NAND2_X1  g542(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n651), .C1(new_n716), .C2(new_n717), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n680), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n645), .A2(new_n464), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n564), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n280), .ZN(G42));
  NOR2_X1   g550(.A1(new_n638), .A2(new_n639), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n650), .A2(new_n418), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT49), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n565), .A2(new_n700), .A3(new_n274), .A4(new_n429), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(new_n630), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n570), .A2(new_n666), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n565), .A2(new_n743), .A3(new_n615), .A4(new_n701), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n733), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT111), .ZN(new_n746));
  INV_X1    g560(.A(new_n738), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n732), .B1(new_n429), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n652), .A2(new_n274), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n744), .A2(new_n630), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT50), .Z(new_n752));
  NAND4_X1  g566(.A1(new_n701), .A2(new_n615), .A3(new_n657), .A4(new_n733), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT112), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n608), .A3(new_n743), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n652), .A2(new_n680), .A3(new_n464), .A4(new_n364), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n737), .A2(new_n574), .A3(new_n584), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n749), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n684), .A2(new_n685), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n754), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT48), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n737), .A2(new_n585), .A3(new_n756), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n652), .A2(new_n275), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n744), .A2(new_n766), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n361), .A2(new_n764), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n759), .A2(new_n760), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n743), .A2(new_n608), .A3(new_n681), .ZN(new_n773));
  INV_X1    g587(.A(new_n357), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n597), .A3(new_n618), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n564), .A2(new_n642), .A3(new_n733), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n698), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n687), .A2(new_n689), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT101), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n777), .B1(new_n781), .B2(new_n686), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n646), .A2(new_n671), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n624), .B2(new_n622), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n676), .A2(new_n651), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n663), .A2(new_n631), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n617), .B(KEYINPUT110), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n459), .A3(new_n607), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n785), .B(new_n789), .C1(new_n638), .C2(new_n639), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n646), .A2(new_n671), .ZN(new_n792));
  AND4_X1   g606(.A1(KEYINPUT52), .A2(new_n625), .A3(new_n792), .A4(new_n790), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n782), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n658), .A2(new_n654), .A3(new_n661), .A4(new_n667), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n695), .A2(new_n653), .B1(new_n564), .B2(new_n660), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n798), .A3(new_n658), .A4(new_n667), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n586), .B1(new_n319), .B2(new_n774), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n276), .A3(new_n587), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n572), .A2(new_n802), .B1(new_n603), .B2(new_n610), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(new_n567), .A3(KEYINPUT109), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT109), .B1(new_n803), .B2(new_n567), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n796), .B(new_n799), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n772), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n777), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n692), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n625), .A2(new_n792), .A3(new_n790), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n784), .A2(KEYINPUT52), .A3(new_n790), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n799), .ZN(new_n815));
  INV_X1    g629(.A(new_n805), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n567), .A3(KEYINPUT109), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n795), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n816), .B2(new_n817), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT54), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n820), .A2(KEYINPUT54), .B1(new_n807), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n771), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(G952), .A2(G953), .ZN(new_n827));
  OAI211_X1 g641(.A(KEYINPUT113), .B(new_n742), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n827), .B1(new_n771), .B2(new_n825), .ZN(new_n830));
  INV_X1    g644(.A(new_n742), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n832), .ZN(G75));
  NOR2_X1   g647(.A1(new_n365), .A2(G952), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT116), .Z(new_n835));
  NAND2_X1  g649(.A1(new_n814), .A2(new_n823), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n353), .B1(new_n807), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(G210), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n263), .B(KEYINPUT114), .Z(new_n840));
  XOR2_X1   g654(.A(new_n266), .B(KEYINPUT55), .Z(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n835), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT56), .B1(new_n838), .B2(KEYINPUT115), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(KEYINPUT115), .B2(new_n838), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n842), .ZN(G51));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT53), .B1(new_n814), .B2(new_n818), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT53), .B(new_n821), .C1(new_n804), .C2(new_n805), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n794), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n794), .A2(new_n851), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n824), .A2(new_n807), .A3(KEYINPUT117), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n424), .B(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(KEYINPUT118), .A3(new_n858), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n648), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n837), .A2(new_n713), .A3(new_n714), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n834), .B1(new_n863), .B2(new_n864), .ZN(G54));
  NAND2_X1  g679(.A1(KEYINPUT58), .A2(G475), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n837), .A2(new_n311), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n311), .B1(new_n837), .B2(new_n867), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n834), .ZN(G60));
  NAND2_X1  g684(.A1(new_n580), .A2(new_n581), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(G478), .A2(G902), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT59), .Z(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n825), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n835), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n874), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n857), .B2(new_n877), .ZN(G63));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT120), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n347), .A2(new_n353), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n880), .B(new_n881), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n807), .B2(new_n836), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n452), .B(KEYINPUT121), .Z(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n606), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n835), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT61), .Z(G66));
  NOR2_X1   g704(.A1(new_n818), .A2(G953), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT122), .ZN(new_n892));
  OAI21_X1  g706(.A(G953), .B1(new_n367), .B2(new_n206), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT123), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n840), .B1(G898), .B2(new_n365), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(G69));
  NAND2_X1  g711(.A1(new_n707), .A2(new_n725), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n762), .A2(new_n786), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n720), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n698), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n735), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n692), .A3(new_n784), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT125), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT125), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n365), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n476), .B1(new_n481), .B2(KEYINPUT30), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n294), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n906), .B(new_n908), .C1(new_n616), .C2(new_n365), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n784), .A2(new_n640), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n911));
  INV_X1    g725(.A(new_n566), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n695), .A2(new_n560), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n430), .A2(new_n800), .A3(new_n627), .A4(new_n733), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n735), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n911), .A2(new_n916), .A3(new_n726), .A4(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT124), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n365), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n909), .B1(new_n920), .B2(new_n908), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n365), .B1(G227), .B2(G900), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n922), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n909), .B(new_n924), .C1(new_n920), .C2(new_n908), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G72));
  NAND2_X1  g740(.A1(G472), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT63), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n544), .A2(new_n525), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n633), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n834), .B1(new_n820), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n904), .A2(new_n818), .A3(new_n905), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n928), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n545), .B(KEYINPUT127), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n928), .B1(new_n919), .B2(new_n806), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT126), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n928), .C1(new_n919), .C2(new_n806), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n525), .B1(new_n482), .B2(new_n485), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(G57));
endmodule


