//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(KEYINPUT64), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(KEYINPUT64), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n221), .A2(G1), .A3(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(G50), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(KEYINPUT1), .B2(new_n218), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  OAI21_X1  g0041(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n242));
  INV_X1    g0042(.A(G150), .ZN(new_n243));
  NOR2_X1   g0043(.A1(G20), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n219), .A2(G33), .A3(new_n220), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  OAI221_X1 g0047(.A(new_n242), .B1(new_n243), .B2(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n249), .A2(new_n253), .A3(new_n250), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n254), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n258), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(G20), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n257), .A2(G50), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n263), .ZN(new_n266));
  INV_X1    g0066(.A(G50), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G274), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(G223), .A3(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(new_n210), .C2(new_n281), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n250), .B1(G33), .B2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n269), .A2(new_n270), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n269), .A2(new_n270), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n287), .A2(G190), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n281), .A2(G232), .A3(G1698), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n286), .ZN(new_n299));
  INV_X1    g0099(.A(new_n276), .ZN(new_n300));
  INV_X1    g0100(.A(new_n279), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(G238), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT13), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n299), .B2(new_n302), .ZN(new_n305));
  OAI21_X1  g0105(.A(G200), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G190), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n244), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n311));
  INV_X1    g0111(.A(G77), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n246), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n255), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n257), .A2(new_n263), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n264), .A2(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n263), .B2(G68), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n266), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n322), .C1(new_n314), .C2(new_n315), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n306), .A2(new_n310), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G169), .B1(new_n304), .B2(new_n305), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT14), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n308), .A2(new_n309), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(G169), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n324), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n269), .B1(new_n287), .B2(G169), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT69), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n287), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n269), .B(KEYINPUT69), .C1(new_n287), .C2(G169), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT70), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n338), .A2(KEYINPUT70), .A3(new_n340), .A4(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT64), .A2(G20), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT64), .A2(G20), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n349), .A2(new_n210), .B1(new_n247), .B2(new_n245), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n246), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n255), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n257), .A2(G77), .A3(new_n263), .A4(new_n264), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n266), .A2(new_n210), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n276), .B1(new_n211), .B2(new_n279), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G107), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n281), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n361), .B2(new_n286), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(G169), .B2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(KEYINPUT71), .B1(new_n339), .B2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n356), .B(new_n365), .C1(G169), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(G190), .ZN(new_n367));
  INV_X1    g0167(.A(new_n362), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n356), .B1(new_n368), .B2(G200), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n364), .A2(new_n366), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n294), .A2(new_n335), .A3(new_n346), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n317), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n247), .B1(new_n258), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n266), .B2(new_n247), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT7), .B1(new_n281), .B2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n349), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(new_n382), .A3(G68), .ZN(new_n383));
  XNOR2_X1  g0183(.A(G58), .B(G68), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(G20), .B1(G159), .B2(new_n244), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n255), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT7), .B1(new_n221), .B2(new_n281), .ZN(new_n390));
  INV_X1    g0190(.A(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n380), .A2(new_n381), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(G68), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n393), .B2(new_n385), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n374), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n275), .A2(G232), .A3(new_n278), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT74), .B1(new_n276), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n276), .A2(new_n397), .A3(KEYINPUT74), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n377), .A2(new_n379), .A3(G226), .A4(G1698), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n377), .A2(new_n379), .A3(G223), .A4(new_n282), .ZN(new_n404));
  INV_X1    g0204(.A(G87), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n404), .C1(new_n376), .C2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(new_n286), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n406), .B2(new_n286), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n401), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(new_n286), .ZN(new_n413));
  AOI21_X1  g0213(.A(G200), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n410), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n406), .A2(new_n407), .A3(new_n286), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n412), .A3(new_n400), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n399), .A3(new_n401), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n288), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT75), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n396), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n415), .B1(new_n410), .B2(new_n414), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(KEYINPUT75), .A3(new_n421), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n395), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT17), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n408), .A2(new_n409), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n411), .A2(G179), .A3(new_n398), .ZN(new_n431));
  INV_X1    g0231(.A(G169), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n430), .A2(new_n431), .B1(new_n432), .B2(new_n420), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n433), .A2(new_n395), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n433), .B2(new_n395), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n425), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n371), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT82), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n377), .A2(new_n379), .A3(G250), .A4(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n377), .A2(new_n379), .A3(G244), .A4(new_n282), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT4), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n444), .A2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n286), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n258), .B(G45), .C1(new_n271), .C2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n454));
  AOI21_X1  g0254(.A(G41), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n450), .B1(new_n455), .B2(KEYINPUT77), .ZN(new_n456));
  AND2_X1   g0256(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT77), .B(new_n271), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G257), .B(new_n275), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n271), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n286), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n464), .A2(new_n466), .A3(new_n459), .A4(new_n450), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n448), .A2(new_n461), .A3(new_n339), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n444), .A2(new_n445), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n442), .A4(new_n443), .ZN(new_n472));
  AOI21_X1  g0272(.A(G179), .B1(new_n472), .B2(new_n286), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n467), .A4(new_n461), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n263), .A2(G97), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n390), .A2(G107), .A3(new_n392), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n245), .A2(new_n312), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n360), .A2(KEYINPUT6), .A3(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n479), .B1(new_n485), .B2(new_n221), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n477), .B1(new_n487), .B2(new_n255), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n258), .A2(G33), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n257), .A2(new_n263), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n448), .A2(new_n461), .A3(new_n467), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n488), .A2(new_n493), .B1(new_n494), .B2(new_n432), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n476), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n448), .A2(new_n461), .A3(G190), .A4(new_n467), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n497), .A2(new_n488), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(G200), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n219), .A2(G33), .A3(G97), .A4(new_n220), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n349), .A2(new_n281), .A3(G68), .ZN(new_n505));
  NAND3_X1  g0305(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n219), .A2(new_n220), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n482), .A2(new_n405), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n255), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n266), .A2(new_n351), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n351), .C2(new_n490), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n258), .A2(G45), .ZN(new_n514));
  INV_X1    g0314(.A(G250), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n275), .C1(G274), .C2(new_n514), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n377), .A2(new_n379), .A3(G238), .A4(new_n282), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n377), .A2(new_n379), .A3(G244), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n281), .A2(new_n523), .A3(G244), .A4(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT80), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n286), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n524), .ZN(new_n528));
  INV_X1    g0328(.A(new_n520), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n528), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n339), .B(new_n517), .C1(new_n527), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n517), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n529), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n275), .B1(new_n533), .B2(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n525), .A2(new_n526), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n513), .B(new_n531), .C1(new_n536), .C2(G169), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n511), .A2(new_n512), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT81), .B1(new_n490), .B2(new_n405), .ZN(new_n539));
  INV_X1    g0339(.A(new_n490), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(G87), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G190), .B(new_n517), .C1(new_n527), .C2(new_n530), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n536), .C2(new_n288), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n441), .B1(new_n501), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n476), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT82), .A3(new_n537), .A4(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n349), .A2(new_n281), .A3(G87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT22), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n349), .A2(new_n281), .A3(new_n552), .A4(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT23), .B1(new_n391), .B2(G107), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G20), .B2(new_n519), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n221), .A2(KEYINPUT85), .A3(new_n558), .A4(new_n360), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n360), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n349), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n557), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n554), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n555), .B1(new_n554), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n255), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n263), .A2(G107), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n540), .B2(G107), .ZN(new_n570));
  OAI211_X1 g0370(.A(G264), .B(new_n275), .C1(new_n456), .C2(new_n460), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n377), .A2(new_n379), .A3(G257), .A4(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n377), .A2(new_n379), .A3(G250), .A4(new_n282), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n286), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n571), .A2(G190), .A3(new_n467), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n467), .A3(new_n576), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n566), .A2(new_n570), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G264), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n581), .B(new_n286), .C1(new_n582), .C2(new_n459), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n576), .A2(new_n467), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n432), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n571), .A2(new_n339), .A3(new_n467), .A4(new_n576), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n566), .B2(new_n570), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n376), .A2(G97), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n219), .A2(new_n590), .A3(new_n220), .A4(new_n443), .ZN(new_n591));
  INV_X1    g0391(.A(G116), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n249), .A2(new_n250), .B1(G20), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n591), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n591), .B2(new_n593), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(G116), .B2(new_n263), .ZN(new_n596));
  AND4_X1   g0396(.A1(G116), .A2(new_n257), .A3(new_n263), .A4(new_n489), .ZN(new_n597));
  OAI21_X1  g0397(.A(G179), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n378), .A2(G33), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n601));
  OAI21_X1  g0401(.A(G303), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n377), .A2(new_n379), .A3(G257), .A4(new_n282), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n377), .A2(new_n379), .A3(G264), .A4(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n599), .B1(new_n605), .B2(new_n286), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n599), .A3(new_n286), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G270), .B(new_n275), .C1(new_n456), .C2(new_n460), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(new_n467), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n598), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n605), .A2(new_n599), .A3(new_n286), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n467), .B(new_n610), .C1(new_n613), .C2(new_n606), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n432), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n596), .B2(new_n597), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n261), .A2(new_n592), .A3(new_n262), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n591), .A2(new_n593), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n591), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n257), .A2(G116), .A3(new_n263), .A4(new_n489), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n432), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n614), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n615), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n619), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT84), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n596), .A2(new_n597), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n614), .B2(new_n400), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n288), .B1(new_n609), .B2(new_n611), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n609), .A2(new_n611), .A3(G190), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n614), .A2(G200), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT84), .A4(new_n632), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n630), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n547), .A2(new_n549), .A3(new_n589), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n440), .A2(new_n640), .ZN(G372));
  NAND2_X1  g0441(.A1(new_n426), .A2(new_n427), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT17), .B1(new_n642), .B2(new_n396), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n424), .B(new_n395), .C1(new_n426), .C2(new_n427), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n332), .B1(new_n327), .B2(KEYINPUT14), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n330), .B1(new_n329), .B2(G169), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n334), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n362), .A2(new_n339), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n366), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n326), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n437), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n294), .B1(new_n344), .B2(new_n345), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n537), .A2(new_n545), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n566), .A2(new_n570), .A3(new_n577), .A4(new_n579), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(KEYINPUT86), .A3(new_n548), .A4(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT86), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n496), .A2(new_n500), .A3(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n546), .ZN(new_n661));
  INV_X1    g0461(.A(new_n630), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n554), .A2(new_n563), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT24), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n554), .A2(new_n563), .A3(new_n555), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n257), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n570), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n586), .B(new_n585), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n658), .A2(new_n661), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n537), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n546), .B2(new_n496), .ZN(new_n673));
  INV_X1    g0473(.A(new_n496), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n537), .A4(new_n545), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n439), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n655), .A2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n258), .A2(G13), .ZN(new_n680));
  OR3_X1    g0480(.A1(new_n221), .A2(KEYINPUT27), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT27), .B1(new_n221), .B2(new_n680), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n632), .ZN(new_n687));
  MUX2_X1   g0487(.A(new_n639), .B(new_n630), .S(new_n687), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n666), .B2(new_n667), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n589), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n668), .B2(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n662), .A2(new_n685), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(new_n589), .B1(new_n588), .B2(new_n686), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n207), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n258), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n508), .A2(G116), .ZN(new_n701));
  INV_X1    g0501(.A(new_n223), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n700), .A2(new_n701), .B1(new_n702), .B2(new_n699), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT87), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n630), .B2(new_n588), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n668), .A2(KEYINPUT89), .A3(new_n629), .A4(new_n619), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n548), .A2(new_n537), .A3(new_n545), .A4(new_n657), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n537), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n673), .A2(new_n675), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT29), .B(new_n686), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n685), .B1(new_n670), .B2(new_n676), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n635), .A2(new_n638), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n589), .A2(new_n662), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n549), .A3(new_n547), .A4(new_n686), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  INV_X1    g0520(.A(new_n494), .ZN(new_n721));
  INV_X1    g0521(.A(new_n578), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n610), .A2(G179), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n609), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n517), .B1(new_n527), .B2(new_n530), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n614), .A2(new_n339), .A3(new_n494), .A4(new_n578), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT88), .B1(new_n728), .B2(new_n536), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n613), .A2(new_n606), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n730), .A2(new_n578), .A3(new_n723), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(KEYINPUT30), .A3(new_n721), .A4(new_n536), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n494), .A2(new_n578), .A3(new_n339), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT88), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n726), .A4(new_n614), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n727), .A2(new_n729), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n685), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n727), .B(new_n732), .C1(new_n536), .C2(new_n728), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n686), .A2(new_n738), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n716), .B1(new_n719), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n715), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n705), .B1(new_n745), .B2(G1), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT90), .Z(G364));
  INV_X1    g0547(.A(G13), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n221), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n700), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n690), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n688), .A2(G330), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT91), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n281), .B(new_n207), .C1(new_n757), .C2(G355), .ZN(new_n758));
  AND2_X1   g0558(.A1(G355), .A2(new_n757), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(G116), .B2(new_n207), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n240), .A2(new_n272), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n698), .A2(new_n281), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n272), .B2(new_n702), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n250), .B1(G20), .B2(new_n432), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n752), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n349), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n773), .A2(new_n339), .A3(G200), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT94), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT94), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n360), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n221), .A2(KEYINPUT93), .A3(G179), .A4(G200), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT93), .ZN(new_n786));
  NAND2_X1  g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n349), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n788), .A3(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n785), .A2(new_n788), .A3(new_n400), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n784), .B1(new_n267), .B2(new_n789), .C1(new_n202), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n774), .A2(G190), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n221), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G97), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n391), .A2(new_n400), .A3(new_n288), .A4(G179), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n281), .B1(new_n800), .B2(new_n405), .ZN(new_n801));
  INV_X1    g0601(.A(new_n210), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n339), .A2(G200), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n773), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n221), .A2(G190), .A3(new_n803), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT92), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n798), .B(new_n805), .C1(new_n201), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n791), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT96), .Z(new_n813));
  INV_X1    g0613(.A(new_n789), .ZN(new_n814));
  INV_X1    g0614(.A(new_n793), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(G326), .B1(G294), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(KEYINPUT97), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n281), .B1(new_n799), .B2(G303), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  INV_X1    g0619(.A(new_n804), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  INV_X1    g0621(.A(G329), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n775), .ZN(new_n823));
  INV_X1    g0623(.A(new_n810), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n819), .B(new_n823), .C1(G322), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n816), .A2(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(new_n782), .ZN(new_n827));
  INV_X1    g0627(.A(new_n790), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n827), .A2(G283), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n813), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n833));
  INV_X1    g0633(.A(new_n769), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n832), .B2(KEYINPUT99), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n772), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT100), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n768), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n688), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n756), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n827), .A2(G87), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n821), .B2(new_n775), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT102), .Z(new_n845));
  NAND2_X1  g0645(.A1(new_n824), .A2(G294), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n380), .B1(new_n800), .B2(new_n360), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n804), .B2(G116), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G283), .A2(new_n828), .B1(new_n814), .B2(G303), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n798), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n281), .B1(new_n800), .B2(new_n267), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G58), .B2(new_n815), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n854), .B2(new_n775), .C1(new_n782), .C2(new_n202), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n824), .A2(G143), .B1(G159), .B2(new_n804), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n857), .B2(new_n789), .C1(new_n243), .C2(new_n790), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(KEYINPUT34), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(KEYINPUT34), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n769), .B1(new_n851), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n769), .A2(new_n766), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n752), .B1(G77), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT103), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n356), .A2(new_n685), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n369), .A2(new_n367), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n651), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(new_n364), .B2(new_n366), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT104), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n651), .A2(new_n870), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n875), .B(new_n876), .C1(new_n370), .C2(new_n870), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n868), .B1(new_n767), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n677), .A2(new_n686), .A3(new_n878), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n714), .B2(new_n878), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(new_n743), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n752), .B1(new_n884), .B2(new_n743), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n881), .A2(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  AOI211_X1 g0688(.A(new_n592), .B(new_n222), .C1(KEYINPUT35), .C2(new_n485), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(KEYINPUT35), .B2(new_n485), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n702), .B1(new_n201), .B2(new_n202), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n892), .A2(new_n210), .B1(G50), .B2(new_n202), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G1), .A3(new_n748), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT106), .Z(new_n896));
  AND2_X1   g0696(.A1(new_n383), .A2(new_n385), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n386), .B(new_n255), .C1(new_n897), .C2(new_n389), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n374), .ZN(new_n899));
  INV_X1    g0699(.A(new_n683), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n438), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n433), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n428), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n683), .B(KEYINPUT107), .Z(new_n908));
  OAI21_X1  g0708(.A(new_n395), .B1(new_n433), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n423), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n395), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n423), .A2(new_n909), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n438), .A2(new_n914), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n912), .B1(KEYINPUT38), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n334), .A2(new_n685), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n648), .A2(new_n325), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n334), .B(new_n685), .C1(new_n333), .C2(new_n326), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n874), .A2(new_n877), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n640), .A2(new_n685), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n737), .A2(new_n738), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n925), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT40), .B1(new_n919), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n921), .A2(new_n922), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n874), .A3(new_n877), .ZN(new_n933));
  INV_X1    g0733(.A(new_n929), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n719), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n901), .B1(new_n645), .B2(new_n437), .ZN(new_n937));
  INV_X1    g0737(.A(new_n911), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n912), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n926), .A2(new_n929), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n440), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n945), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n946), .A2(new_n947), .A3(new_n716), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n651), .A2(new_n685), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n883), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n940), .A3(new_n932), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n903), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n438), .A2(new_n914), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n916), .A2(new_n910), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n333), .A2(new_n334), .A3(new_n686), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n437), .A2(new_n908), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n952), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n713), .B(new_n439), .C1(KEYINPUT29), .C2(new_n714), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n655), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n948), .A2(new_n967), .B1(new_n258), .B2(new_n749), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n948), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n896), .B1(new_n968), .B2(new_n969), .ZN(G367));
  NAND2_X1  g0770(.A1(new_n233), .A2(new_n762), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n770), .C1(new_n207), .C2(new_n351), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n752), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n543), .A2(new_n686), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n671), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n546), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n839), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n775), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n800), .A2(new_n592), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n380), .B1(new_n360), .B2(new_n793), .C1(new_n980), .C2(KEYINPUT46), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n981), .C1(G283), .C2(new_n804), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT109), .Z(new_n984));
  INV_X1    g0784(.A(G303), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n982), .B(new_n984), .C1(new_n985), .C2(new_n810), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n782), .A2(new_n491), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G311), .B2(new_n814), .ZN(new_n988));
  INV_X1    g0788(.A(G294), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n790), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n796), .A2(new_n202), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G150), .B2(new_n824), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n281), .B1(new_n800), .B2(new_n201), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n804), .B2(G50), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(new_n857), .C2(new_n775), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n827), .A2(new_n802), .B1(G143), .B2(new_n814), .ZN(new_n996));
  INV_X1    g0796(.A(G159), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n790), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n986), .A2(new_n990), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n973), .B(new_n977), .C1(new_n1000), .C2(new_n769), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n750), .A2(G1), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n686), .B1(new_n493), .B2(new_n488), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n501), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n496), .A2(new_n686), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n696), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT45), .Z(new_n1010));
  NOR2_X1   g0810(.A1(new_n1008), .A2(new_n696), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT44), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n694), .C2(KEYINPUT108), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n694), .A2(KEYINPUT108), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n695), .A2(new_n589), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n693), .B2(new_n695), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n689), .B(new_n1017), .Z(new_n1018));
  AOI21_X1  g0818(.A(new_n744), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n699), .B(KEYINPUT41), .Z(new_n1020));
  OAI21_X1  g0820(.A(new_n1003), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n588), .A2(new_n500), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n685), .B1(new_n1024), .B2(new_n496), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1022), .B2(KEYINPUT42), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1023), .A2(new_n1026), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n694), .A2(new_n1007), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1029), .B(new_n1030), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n1001), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(G387));
  AOI21_X1  g0833(.A(new_n763), .B1(new_n230), .B2(G45), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n701), .B(new_n272), .C1(new_n202), .C2(new_n312), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(KEYINPUT110), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n247), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(KEYINPUT110), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1034), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n281), .A2(new_n207), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1042), .B1(G107), .B2(new_n207), .C1(new_n701), .C2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n751), .B1(new_n1044), .B2(new_n770), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n693), .B2(new_n839), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n790), .A2(new_n247), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1047), .B(new_n987), .C1(G159), .C2(new_n814), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n799), .A2(new_n802), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n281), .B(new_n1049), .C1(new_n775), .C2(new_n243), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G68), .B2(new_n804), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n796), .A2(new_n351), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n824), .B2(G50), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n281), .B1(new_n776), .B2(G326), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n824), .A2(G317), .B1(G303), .B2(new_n804), .ZN(new_n1056));
  INV_X1    g0856(.A(G322), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n821), .A2(new_n790), .B1(new_n789), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n815), .A2(G283), .B1(G294), .B2(new_n799), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1055), .B1(new_n592), .B2(new_n782), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1054), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1046), .B1(new_n1070), .B2(new_n769), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT113), .Z(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1002), .B2(new_n1018), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n745), .A2(new_n1018), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n745), .A2(new_n1018), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n699), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(new_n699), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1075), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1015), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1079), .B2(new_n1015), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n281), .B1(new_n799), .B2(G283), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n793), .B2(new_n592), .C1(new_n775), .C2(new_n1057), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1084), .B(new_n783), .C1(G294), .C2(new_n804), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n810), .A2(new_n821), .B1(new_n978), .B2(new_n789), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n985), .C2(new_n790), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n810), .A2(new_n997), .B1(new_n243), .B2(new_n789), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n796), .A2(new_n312), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n281), .B1(new_n202), .B2(new_n800), .C1(new_n820), .C2(new_n247), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G143), .C2(new_n776), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n828), .A2(G50), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1090), .A2(new_n1093), .A3(new_n843), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n834), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n237), .A2(new_n762), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n771), .B1(G97), .B2(new_n698), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n751), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT114), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n768), .B2(new_n1007), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1015), .B2(new_n1002), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1081), .A2(new_n1082), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1082), .B1(new_n1081), .B2(new_n1102), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  NAND3_X1  g0907(.A1(new_n874), .A2(new_n686), .A3(new_n877), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n670), .B2(new_n676), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n932), .B1(new_n1109), .B2(new_n949), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n960), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n958), .A2(new_n959), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n878), .B(new_n686), .C1(new_n711), .C2(new_n712), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n923), .B1(new_n1114), .B2(new_n950), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n960), .B1(new_n954), .B2(new_n957), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n742), .A2(new_n878), .A3(new_n932), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1113), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n960), .A2(new_n1110), .B1(new_n958), .B2(new_n959), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n925), .B(G330), .C1(new_n926), .C2(new_n929), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1002), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1120), .A2(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1002), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(G330), .B(new_n439), .C1(new_n926), .C2(new_n929), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n713), .A2(new_n439), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT29), .B1(new_n677), .B2(new_n686), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n655), .B(new_n1135), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n965), .A2(KEYINPUT117), .A3(new_n655), .A4(new_n1135), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1114), .A2(new_n950), .ZN(new_n1143));
  OAI211_X1 g0943(.A(G330), .B(new_n878), .C1(new_n926), .C2(new_n929), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n923), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n716), .B(new_n924), .C1(new_n719), .C2(new_n741), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1126), .B1(new_n1146), .B2(new_n932), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1145), .A2(new_n1119), .B1(new_n1147), .B2(new_n951), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT118), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n951), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1144), .A2(new_n923), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n950), .A3(new_n1114), .A4(new_n1119), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n699), .B(new_n1150), .C1(new_n1158), .C2(new_n1132), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1112), .A2(new_n766), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n863), .A2(new_n247), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n827), .A2(G50), .B1(G137), .B2(new_n828), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n789), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n824), .A2(G132), .B1(new_n797), .B2(G159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n380), .B1(new_n776), .B2(G125), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT53), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n800), .B2(new_n243), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n799), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1168), .A2(new_n1169), .B1(new_n804), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1164), .A2(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT120), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT120), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n281), .B1(new_n799), .B2(G87), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n989), .B2(new_n775), .C1(new_n820), .C2(new_n491), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1091), .B(new_n1178), .C1(G116), .C2(new_n824), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n827), .A2(G68), .B1(G283), .B2(new_n814), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n360), .C2(new_n790), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1176), .A3(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n751), .B(new_n1161), .C1(new_n1182), .C2(new_n769), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1160), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1134), .A2(new_n1159), .A3(new_n1184), .ZN(G378));
  NAND2_X1  g0985(.A1(new_n294), .A2(new_n342), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n269), .A2(new_n900), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT122), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n767), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n790), .A2(new_n854), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n804), .A2(G137), .B1(new_n799), .B2(new_n1171), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n796), .B2(new_n243), .C1(new_n810), .C2(new_n1163), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G125), .C2(new_n814), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n827), .A2(G159), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n376), .A2(new_n271), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n776), .B2(G124), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n827), .A2(G58), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n491), .B2(new_n790), .C1(new_n592), .C2(new_n789), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n824), .A2(G107), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n776), .A2(G283), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n281), .A2(G41), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1049), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(new_n351), .C2(new_n820), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1206), .A2(new_n1208), .A3(new_n991), .A4(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n267), .B(new_n1202), .C1(new_n281), .C2(G41), .ZN(new_n1216));
  AND4_X1   g1016(.A1(new_n1204), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n752), .B1(G50), .B2(new_n864), .C1(new_n1217), .C2(new_n834), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1193), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n941), .B1(new_n935), .B2(new_n918), .ZN(new_n1221));
  OAI21_X1  g1021(.A(G330), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n964), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n716), .B1(new_n931), .B2(new_n942), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n952), .A2(new_n962), .A3(new_n963), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1226), .A3(new_n1192), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1192), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1219), .B1(new_n1230), .B2(new_n1002), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1150), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1190), .B(new_n1191), .Z(new_n1235));
  NOR2_X1   g1035(.A1(new_n964), .A2(new_n1222), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(KEYINPUT57), .A3(new_n1227), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1142), .B1(new_n1132), .B2(new_n1149), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n699), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1231), .B1(new_n1234), .B2(new_n1241), .ZN(G375));
  OAI21_X1  g1042(.A(new_n752), .B1(G68), .B2(new_n864), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n281), .B1(new_n799), .B2(G97), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n985), .B2(new_n775), .C1(new_n820), .C2(new_n360), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1052), .B(new_n1245), .C1(G283), .C2(new_n824), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G116), .A2(new_n828), .B1(new_n814), .B2(G294), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(new_n312), .C2(new_n782), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n824), .A2(G137), .B1(new_n828), .B2(new_n1171), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n854), .B2(new_n789), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n797), .A2(G50), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n804), .A2(G150), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n281), .B1(new_n800), .B2(new_n997), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n776), .B2(G128), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1205), .A2(new_n1252), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1248), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1243), .B1(new_n1257), .B2(new_n769), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n767), .B2(new_n932), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1148), .B2(new_n1003), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1020), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1158), .B2(new_n1264), .ZN(G381));
  OR2_X1    g1065(.A1(G396), .A2(G393), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G384), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1106), .A2(new_n1032), .A3(new_n1267), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G378), .A2(new_n1268), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1069(.A(G378), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n684), .A2(G213), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  XNOR2_X1  g1073(.A(new_n841), .B(G393), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT126), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1032), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1105), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G387), .A2(new_n1277), .A3(new_n1103), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1278), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1276), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1274), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1231), .C1(new_n1234), .C2(new_n1241), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1151), .A3(new_n1157), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1078), .B1(new_n1132), .B2(new_n1149), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1289), .A2(new_n1290), .B1(new_n1160), .B2(new_n1183), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1238), .A2(new_n1227), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1292), .A2(new_n1240), .A3(new_n1020), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1292), .A2(new_n1003), .B1(new_n1193), .B2(new_n1218), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1134), .B(new_n1291), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1271), .B1(new_n1287), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1078), .B1(new_n1232), .B2(new_n1155), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1262), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1142), .A2(new_n1148), .A3(KEYINPUT60), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1297), .A2(new_n1299), .A3(new_n1303), .A4(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1305), .B2(new_n1261), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n887), .B(new_n1260), .C1(new_n1302), .C2(new_n1304), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n699), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1303), .B1(new_n1312), .B2(new_n1300), .ZN(new_n1313));
  AND4_X1   g1113(.A1(new_n1303), .A2(new_n1297), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1261), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n887), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(G384), .A3(new_n1261), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1296), .B1(new_n1309), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1296), .B(new_n1321), .C1(new_n1309), .C2(new_n1318), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1271), .A2(G2897), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1287), .A2(new_n1295), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1328), .B2(new_n1271), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1308), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1316), .A2(KEYINPUT125), .A3(new_n1317), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1326), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1329), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1286), .B1(new_n1323), .B2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1285), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1282), .B2(new_n1275), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1325), .B1(new_n1309), .B2(new_n1318), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1325), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1296), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT61), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1319), .A2(new_n1341), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1296), .B(KEYINPUT63), .C1(new_n1309), .C2(new_n1318), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1336), .A2(new_n1340), .A3(new_n1342), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1334), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1270), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1287), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1348));
  OR3_X1    g1148(.A1(new_n1347), .A2(KEYINPUT127), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT127), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1350));
  AOI22_X1  g1150(.A1(new_n1330), .A2(new_n1331), .B1(new_n1346), .B2(new_n1287), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1336), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1286), .B(new_n1349), .C1(new_n1351), .C2(new_n1350), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


