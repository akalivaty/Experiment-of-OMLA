//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  AOI21_X1  g000(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT97), .ZN(new_n204));
  XNOR2_X1  g003(.A(G99gat), .B(G106gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206));
  INV_X1    g005(.A(G85gat), .ZN(new_n207));
  INV_X1    g006(.A(G92gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(KEYINPUT8), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(G85gat), .A3(G92gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(new_n204), .B(new_n205), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n209), .ZN(new_n217));
  INV_X1    g016(.A(new_n205), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n209), .A3(new_n205), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n204), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G50gat), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G43gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(G43gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(G50gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT84), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(KEYINPUT15), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT85), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G36gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n238), .A3(G29gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT14), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  INV_X1    g040(.A(G29gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n235), .A3(KEYINPUT14), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(KEYINPUT86), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n234), .B(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n227), .A2(new_n229), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT87), .B(KEYINPUT15), .Z(new_n248));
  NOR3_X1   g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n223), .B(new_n224), .C1(new_n245), .C2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n251), .A3(KEYINPUT86), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n244), .A2(KEYINPUT15), .A3(new_n233), .A4(new_n230), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT88), .A2(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n223), .A2(new_n224), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n222), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n254), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n214), .A2(new_n205), .A3(new_n209), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n205), .B1(new_n214), .B2(new_n209), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n215), .B1(new_n262), .B2(new_n204), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G190gat), .B(G218gat), .Z(new_n268));
  OAI21_X1  g067(.A(KEYINPUT99), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n253), .ZN(new_n270));
  INV_X1    g069(.A(new_n249), .ZN(new_n271));
  AND4_X1   g070(.A1(new_n270), .A2(new_n271), .A3(new_n255), .A4(new_n256), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n256), .B1(new_n254), .B2(new_n255), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n264), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n265), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT99), .ZN(new_n277));
  INV_X1    g076(.A(new_n268), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G134gat), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n274), .A2(new_n268), .A3(new_n275), .A4(new_n265), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n258), .A2(new_n266), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(KEYINPUT98), .A3(new_n268), .A4(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n280), .A2(new_n281), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n280), .B2(new_n287), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT96), .B(G162gat), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n267), .A2(KEYINPUT99), .A3(new_n268), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n284), .A2(new_n286), .ZN(new_n296));
  OAI21_X1  g095(.A(G134gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n287), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n203), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n292), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n202), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G71gat), .ZN(new_n305));
  INV_X1    g104(.A(G78gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G71gat), .A2(G78gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G57gat), .B(G64gat), .Z(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(KEYINPUT9), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT92), .ZN(new_n312));
  INV_X1    g111(.A(G57gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n312), .B(G64gat), .C1(new_n313), .C2(KEYINPUT93), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n315));
  INV_X1    g114(.A(G64gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n315), .B(G57gat), .C1(new_n316), .C2(KEYINPUT92), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT92), .B1(new_n316), .B2(G57gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT9), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n308), .B1(new_n307), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT94), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(KEYINPUT94), .A3(new_n321), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT21), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT89), .ZN(new_n329));
  XNOR2_X1  g128(.A(G15gat), .B(G22gat), .ZN(new_n330));
  INV_X1    g129(.A(G1gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT16), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n330), .A2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n329), .B(G8gat), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(G8gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n329), .A2(G8gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(new_n332), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n335), .A2(KEYINPUT91), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT91), .B1(new_n335), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(KEYINPUT21), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G155gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n344), .B(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(G231gat), .A2(G233gat), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n328), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n328), .A3(new_n350), .ZN(new_n353));
  XNOR2_X1  g152(.A(G183gat), .B(G211gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT20), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n352), .B2(new_n353), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n304), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G230gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT97), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT10), .B1(new_n364), .B2(new_n215), .ZN(new_n365));
  INV_X1    g164(.A(new_n311), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n319), .A2(KEYINPUT94), .A3(new_n321), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT94), .B1(new_n319), .B2(new_n321), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n326), .A2(new_n222), .A3(KEYINPUT100), .A4(KEYINPUT10), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n222), .A2(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n219), .A2(new_n220), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(new_n366), .C1(new_n368), .C2(new_n367), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT10), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n362), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT102), .ZN(new_n378));
  INV_X1    g177(.A(new_n362), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT102), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n362), .C1(new_n372), .C2(new_n376), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G120gat), .B(G148gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT101), .ZN(new_n385));
  INV_X1    g184(.A(G176gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G204gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n377), .A2(new_n380), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G141gat), .B(G148gat), .Z(new_n394));
  INV_X1    g193(.A(G155gat), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT2), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G155gat), .B(G162gat), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n398), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G197gat), .B(G204gat), .ZN(new_n406));
  INV_X1    g205(.A(G211gat), .ZN(new_n407));
  INV_X1    g206(.A(G218gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(KEYINPUT22), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n398), .B(new_n399), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n402), .B1(new_n412), .B2(KEYINPUT29), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n405), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(G22gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT31), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(new_n228), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  OR3_X1    g222(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(KEYINPUT78), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G226gat), .ZN(new_n428));
  INV_X1    g227(.A(G233gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT27), .B(G183gat), .ZN(new_n433));
  INV_X1    g232(.A(G190gat), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g235(.A(G169gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(new_n386), .ZN(new_n438));
  NOR2_X1   g237(.A1(G169gat), .A2(G176gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(KEYINPUT26), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n439), .B(KEYINPUT66), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT26), .ZN(new_n443));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n436), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n439), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT23), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n438), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(KEYINPUT24), .ZN(new_n452));
  NOR2_X1   g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n444), .A2(KEYINPUT24), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n449), .A2(KEYINPUT25), .A3(new_n451), .A4(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n440), .ZN(new_n459));
  INV_X1    g258(.A(new_n438), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n444), .A2(KEYINPUT24), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n439), .A2(KEYINPUT23), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n462), .B(new_n463), .C1(new_n453), .C2(new_n452), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n458), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n431), .B1(new_n446), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n404), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n470), .A2(KEYINPUT73), .A3(new_n431), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT73), .B1(new_n470), .B2(new_n431), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n412), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n470), .B2(new_n431), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(new_n412), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT74), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(KEYINPUT74), .A3(new_n475), .ZN(new_n479));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(new_n316), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(new_n208), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT75), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n476), .A2(KEYINPUT75), .A3(KEYINPUT30), .A4(new_n484), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n491));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT0), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G57gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(new_n207), .ZN(new_n495));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G113gat), .B(G120gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G127gat), .B(G134gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT1), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT1), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT69), .B(G120gat), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n505), .A2(G113gat), .ZN(new_n506));
  INV_X1    g305(.A(G113gat), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(G120gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n502), .B(new_n503), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n501), .B1(new_n509), .B2(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n401), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n413), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n497), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n413), .A2(KEYINPUT3), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n403), .A3(new_n511), .A4(new_n512), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT4), .B(new_n413), .C1(new_n511), .C2(new_n512), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(new_n496), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT5), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n495), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n524), .A2(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(new_n495), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533));
  OAI211_X1 g332(.A(KEYINPUT77), .B(new_n495), .C1(new_n524), .C2(new_n526), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n529), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n531), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n490), .A2(new_n491), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT30), .B1(new_n476), .B2(new_n484), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n489), .B2(KEYINPUT76), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n427), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n469), .A2(new_n513), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n511), .A2(new_n446), .A3(new_n466), .A4(new_n512), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n541), .A2(G227gat), .A3(G233gat), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT32), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G43gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G71gat), .ZN(new_n549));
  INV_X1    g348(.A(G99gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n551), .A2(KEYINPUT33), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT71), .B1(new_n544), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n542), .ZN(new_n557));
  INV_X1    g356(.A(G227gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n429), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT34), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(KEYINPUT71), .C1(new_n544), .C2(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n560), .A3(new_n552), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT72), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n556), .A2(new_n561), .A3(KEYINPUT72), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT36), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT79), .B1(new_n540), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n535), .A2(new_n536), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n483), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n539), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n427), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578));
  INV_X1    g377(.A(new_n571), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n474), .A2(new_n412), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n471), .A2(new_n472), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n467), .ZN(new_n583));
  OAI211_X1 g382(.A(KEYINPUT37), .B(new_n581), .C1(new_n583), .C2(new_n412), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n476), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n482), .A4(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n535), .A2(new_n536), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n478), .A2(KEYINPUT37), .A3(new_n479), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n482), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT38), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n476), .A2(new_n484), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(KEYINPUT38), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n589), .A2(new_n593), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n538), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n483), .A2(new_n487), .A3(new_n598), .A4(new_n488), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n497), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n601), .A2(KEYINPUT39), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n514), .A2(new_n515), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(KEYINPUT39), .C1(new_n497), .C2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n604), .A3(new_n495), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT40), .A4(new_n495), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n608), .A2(new_n532), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n599), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n610), .A2(new_n427), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n597), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n572), .A2(new_n580), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n566), .A2(new_n567), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n427), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT35), .B1(new_n575), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n599), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT35), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n617), .A2(new_n573), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT81), .ZN(new_n620));
  INV_X1    g419(.A(new_n565), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n560), .B1(new_n564), .B2(new_n552), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT81), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(new_n427), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n616), .A2(new_n626), .ZN(new_n627));
  AOI211_X1 g426(.A(new_n361), .B(new_n393), .C1(new_n613), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n250), .A2(new_n257), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n335), .A2(new_n339), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n340), .A2(new_n341), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n254), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT90), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n629), .A2(new_n630), .B1(new_n632), .B2(new_n254), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n342), .A2(new_n259), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n635), .B(KEYINPUT13), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT82), .B(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT11), .B(G169gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n640), .A3(new_n652), .A4(new_n644), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n573), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n331), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n617), .ZN(new_n660));
  NOR2_X1   g459(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n660), .A2(new_n666), .A3(new_n662), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n657), .B2(new_n617), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1325gat));
  AND2_X1   g470(.A1(new_n628), .A2(new_n656), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n623), .A2(new_n624), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(G15gat), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n571), .A2(G15gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT104), .Z(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n672), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n657), .A2(new_n427), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  AOI21_X1  g480(.A(new_n304), .B1(new_n613), .B2(new_n627), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n360), .A2(new_n393), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n656), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n573), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n242), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n613), .A2(new_n627), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n301), .A2(new_n302), .A3(new_n202), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n202), .B1(new_n301), .B2(new_n302), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(KEYINPUT44), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n612), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n627), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n692), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n656), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n655), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n693), .A2(new_n683), .A3(new_n699), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n573), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n706), .ZN(G1328gat));
  NAND2_X1  g506(.A1(new_n236), .A2(new_n238), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n684), .A2(new_n709), .A3(new_n617), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n712), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n705), .B2(new_n617), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n571), .A2(G43gat), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n226), .B1(new_n684), .B2(new_n673), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT47), .B1(new_n718), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n705), .B2(new_n427), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n576), .A2(new_n228), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n685), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n393), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n695), .B2(new_n627), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n361), .A2(new_n704), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n573), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n313), .ZN(G1332gat));
  AND2_X1   g535(.A1(new_n732), .A2(new_n733), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n599), .B(KEYINPUT108), .Z(new_n738));
  AND2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g542(.A1(new_n737), .A2(G71gat), .A3(new_n571), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n305), .B1(new_n734), .B2(new_n673), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT109), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n427), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(new_n306), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n360), .A2(new_n704), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n696), .A2(new_n692), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n696), .A2(new_n755), .A3(KEYINPUT51), .A4(new_n692), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n686), .A3(new_n393), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n360), .A2(new_n704), .A3(new_n731), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n693), .A2(new_n699), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n573), .A2(new_n207), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n761), .A2(new_n207), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n760), .A2(new_n208), .A3(new_n393), .A4(new_n738), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n763), .A2(new_n738), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n208), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n693), .A2(new_n599), .A3(new_n699), .A4(new_n762), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n767), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n772), .B2(KEYINPUT52), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n774), .B(new_n766), .C1(new_n771), .C2(new_n767), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n773), .B2(new_n775), .ZN(G1337gat));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n393), .A3(new_n674), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n579), .A2(new_n550), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(new_n550), .B1(new_n763), .B2(new_n778), .ZN(G1338gat));
  NAND4_X1  g578(.A1(new_n693), .A2(new_n576), .A3(new_n699), .A4(new_n762), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n427), .A2(G106gat), .A3(new_n731), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT111), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n780), .A2(G106gat), .B1(new_n760), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT53), .Z(G1339gat));
  NAND4_X1  g583(.A1(new_n304), .A2(new_n360), .A3(new_n731), .A4(new_n703), .ZN(new_n785));
  INV_X1    g584(.A(new_n392), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT54), .B1(new_n378), .B2(new_n382), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n375), .B1(new_n263), .B2(new_n326), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT10), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n370), .A3(new_n371), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT54), .B1(new_n791), .B2(new_n362), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n370), .A2(new_n371), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n379), .B1(new_n793), .B2(new_n790), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n389), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT55), .B1(new_n787), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n372), .A2(new_n376), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n379), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n391), .B1(new_n799), .B2(new_n377), .ZN(new_n800));
  INV_X1    g599(.A(new_n382), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n381), .B1(new_n791), .B2(new_n362), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n786), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n639), .A2(new_n635), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n642), .A2(new_n643), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n650), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT112), .B(new_n650), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n655), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n300), .A2(new_n303), .A3(new_n806), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n701), .A2(new_n806), .A3(new_n702), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n393), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n690), .B2(new_n691), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n785), .B1(new_n820), .B2(new_n360), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n738), .A2(new_n573), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n625), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n656), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n615), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n826), .A3(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n704), .A2(new_n507), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT113), .ZN(G1340gat));
  OAI21_X1  g629(.A(G120gat), .B1(new_n823), .B2(new_n731), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n393), .A2(new_n505), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n827), .B2(new_n832), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834));
  INV_X1    g633(.A(new_n360), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n823), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n827), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n360), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n834), .B2(new_n838), .ZN(G1342gat));
  OAI21_X1  g638(.A(G134gat), .B1(new_n823), .B2(new_n304), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n821), .A2(new_n617), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n304), .A2(new_n573), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n281), .A3(new_n826), .A4(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n738), .A2(new_n573), .A3(new_n571), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n813), .A2(new_n731), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n787), .A2(new_n795), .A3(KEYINPUT55), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n804), .B1(new_n800), .B2(new_n803), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n392), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n824), .B1(new_n856), .B2(KEYINPUT116), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n806), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n853), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT117), .B1(new_n692), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n859), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n656), .B1(new_n806), .B2(new_n858), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n817), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n304), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n861), .A2(new_n815), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n835), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n852), .B1(new_n868), .B2(new_n785), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n821), .B2(new_n576), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n704), .B(new_n851), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n821), .A2(new_n576), .ZN(new_n874));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n656), .A4(new_n851), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n850), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n850), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n656), .B(new_n851), .C1(new_n869), .C2(new_n871), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(G141gat), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT118), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(G141gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n821), .A2(new_n576), .A3(new_n851), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G141gat), .A3(new_n824), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n872), .B2(G141gat), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n886), .B(new_n887), .C1(new_n850), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n881), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n851), .B1(new_n869), .B2(new_n871), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n891), .B(G148gat), .C1(new_n892), .C2(new_n731), .ZN(new_n893));
  INV_X1    g692(.A(new_n785), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n360), .B1(new_n815), .B2(new_n819), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n576), .B(new_n870), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n815), .B1(new_n692), .B2(new_n860), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n835), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n304), .A2(new_n824), .A3(new_n360), .A4(new_n731), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n427), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n851), .B(KEYINPUT119), .Z(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n393), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n904), .B2(KEYINPUT59), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  AOI211_X1 g705(.A(new_n906), .B(new_n891), .C1(new_n903), .C2(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n893), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n883), .A2(G148gat), .A3(new_n731), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1345gat));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n395), .A3(new_n835), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n874), .A2(new_n360), .A3(new_n851), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n395), .B2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n892), .B2(new_n304), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n579), .A2(new_n576), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n841), .A2(new_n396), .A3(new_n842), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n686), .A2(new_n617), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT121), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(KEYINPUT121), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n821), .A2(new_n625), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n824), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n821), .A2(new_n573), .A3(new_n826), .A4(new_n738), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n704), .A2(new_n437), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G1348gat));
  NOR3_X1   g725(.A1(new_n922), .A2(new_n386), .A3(new_n731), .ZN(new_n927));
  INV_X1    g726(.A(new_n924), .ZN(new_n928));
  AOI21_X1  g727(.A(G176gat), .B1(new_n928), .B2(new_n393), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1349gat));
  OR3_X1    g731(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n835), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n922), .B2(new_n835), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(G183gat), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n433), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT123), .A3(new_n360), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT123), .B1(new_n937), .B2(new_n360), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n935), .B(new_n942), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n922), .B2(new_n304), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n434), .A3(new_n692), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n821), .A2(new_n738), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n686), .A3(new_n915), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n704), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n919), .A2(new_n920), .A3(new_n571), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n901), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n656), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n950), .A2(new_n388), .A3(new_n393), .A4(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n901), .A2(new_n393), .A3(new_n953), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n961), .B(new_n962), .C1(new_n388), .C2(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n950), .A2(new_n407), .A3(new_n360), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT126), .Z(new_n966));
  NAND3_X1  g765(.A1(new_n901), .A2(new_n360), .A3(new_n953), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n901), .A2(new_n969), .A3(new_n360), .A4(new_n953), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(G211gat), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT63), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n968), .A2(new_n973), .A3(G211gat), .A4(new_n970), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n966), .A2(new_n972), .A3(new_n974), .ZN(G1354gat));
  AOI21_X1  g774(.A(G218gat), .B1(new_n950), .B2(new_n692), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n304), .A2(new_n408), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n954), .B2(new_n977), .ZN(G1355gat));
endmodule


