//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n188), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT66), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G137), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G134), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n201), .A2(G134), .B1(G137), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT64), .A2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT64), .A2(G134), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n205), .A2(new_n206), .A3(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n207), .B2(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(new_n206), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT64), .A2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n197), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT65), .A3(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n203), .A2(new_n208), .A3(new_n215), .A4(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(G116), .B(G119), .Z(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n219), .A3(new_n221), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n218), .A3(G143), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n220), .B(G146), .C1(new_n238), .C2(KEYINPUT1), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n198), .A2(new_n200), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n215), .B1(new_n211), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT67), .B1(new_n216), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n229), .A2(new_n237), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n227), .B1(new_n214), .B2(new_n216), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n216), .A2(new_n247), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT30), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n229), .A2(new_n249), .A3(new_n250), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(KEYINPUT30), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n195), .B(new_n251), .C1(new_n257), .C2(new_n237), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n261));
  NOR4_X1   g075(.A1(new_n252), .A2(new_n261), .A3(new_n248), .A4(new_n236), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n229), .A2(new_n263), .A3(new_n253), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n252), .A2(new_n261), .A3(new_n248), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(new_n263), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n266), .B2(new_n236), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n195), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n237), .B1(new_n229), .B2(new_n253), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT28), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n252), .A2(new_n254), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT28), .B1(new_n274), .B2(new_n237), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n236), .B1(new_n252), .B2(new_n254), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n251), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n194), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(G472), .A2(G902), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT32), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  INV_X1    g100(.A(new_n284), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n286), .B(new_n287), .C1(new_n269), .C2(new_n282), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n187), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n260), .A2(new_n268), .B1(new_n281), .B2(new_n194), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n281), .B2(new_n194), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n272), .B(new_n277), .C1(new_n251), .C2(new_n278), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT71), .A3(new_n195), .A4(new_n276), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  INV_X1    g113(.A(new_n267), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n194), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n294), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n256), .A2(new_n236), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n251), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n275), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n194), .A2(new_n299), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G472), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n289), .A2(new_n292), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G140), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G125), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(KEYINPUT73), .A3(G140), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(G125), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n320), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(new_n218), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n311), .A2(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n325), .A3(new_n218), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n328), .B(KEYINPUT72), .Z(new_n329));
  NOR2_X1   g143(.A1(new_n238), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G119), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G128), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n329), .B(new_n331), .C1(KEYINPUT23), .C2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n330), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT24), .B(G110), .Z(new_n336));
  OAI22_X1  g150(.A1(new_n334), .A2(G110), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n323), .B(new_n218), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n334), .A2(G110), .B1(new_n335), .B2(new_n336), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n327), .A2(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT75), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT25), .B1(new_n347), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  INV_X1    g163(.A(G902), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(G234), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n345), .A2(new_n352), .A3(new_n350), .A4(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT76), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n347), .A2(KEYINPUT76), .A3(new_n356), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G952), .ZN(new_n360));
  AOI211_X1 g174(.A(G953), .B(new_n360), .C1(G234), .C2(G237), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n350), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT21), .B(G898), .Z(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G469), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n190), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT77), .B1(new_n371), .B2(G104), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n374), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n371), .A3(G104), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n383), .A3(G101), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n377), .A2(new_n379), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n376), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n385), .B2(new_n376), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(new_n383), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n389), .B2(new_n383), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .A4(new_n387), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n227), .B(new_n382), .C1(new_n391), .C2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n374), .A2(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n371), .A2(G104), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n243), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n403), .B(KEYINPUT10), .Z(new_n404));
  OAI21_X1  g218(.A(new_n217), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(new_n396), .ZN(new_n406));
  INV_X1    g220(.A(new_n382), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n228), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n403), .B(KEYINPUT10), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n214), .A2(new_n410), .A3(new_n216), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n214), .B2(new_n216), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n370), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n387), .A2(new_n400), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n243), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n403), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n217), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n414), .A2(new_n370), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n367), .B(new_n350), .C1(new_n415), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n414), .A2(new_n423), .ZN(new_n426));
  INV_X1    g240(.A(new_n370), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n405), .A2(new_n414), .A3(new_n370), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(G469), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(G469), .A2(G902), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT9), .B(G234), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G221), .B1(new_n435), .B2(G902), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G214), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n438), .A2(G237), .A3(G953), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(G143), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT85), .B(G143), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n441), .B(new_n215), .C1(new_n439), .C2(new_n442), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT86), .A3(new_n445), .ZN(new_n446));
  OR3_X1    g260(.A1(new_n443), .A2(KEYINPUT86), .A3(G131), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT17), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(KEYINPUT17), .A3(G131), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT88), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n448), .A2(new_n450), .A3(new_n338), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n374), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n443), .A2(KEYINPUT18), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n326), .B1(new_n317), .B2(new_n218), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n443), .A2(KEYINPUT18), .A3(G131), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n455), .A2(new_n445), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n451), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n447), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT19), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n320), .A2(new_n325), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n317), .B2(new_n464), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n466), .A2(G146), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT87), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n463), .A2(new_n324), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n453), .B1(new_n469), .B2(new_n458), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT89), .Z(new_n473));
  OAI21_X1  g287(.A(KEYINPUT20), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n475));
  INV_X1    g289(.A(new_n473), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(new_n476), .C1(new_n460), .C2(new_n470), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n451), .A2(new_n459), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n453), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n350), .B1(new_n480), .B2(new_n460), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G475), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT13), .B1(new_n220), .B2(G128), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT90), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n220), .A2(G128), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n220), .A2(G128), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G134), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n202), .ZN(new_n493));
  XNOR2_X1  g307(.A(G116), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n371), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n496), .A2(KEYINPUT91), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G122), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G116), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n371), .B1(new_n501), .B2(KEYINPUT14), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n499), .A2(new_n502), .B1(new_n371), .B2(new_n494), .ZN(new_n503));
  INV_X1    g317(.A(new_n493), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n492), .A2(new_n202), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n496), .A2(KEYINPUT91), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n435), .A2(new_n349), .A3(G953), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n497), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n513), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n513), .B(KEYINPUT92), .C1(KEYINPUT15), .C2(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n483), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT83), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT5), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n332), .A3(G116), .ZN(new_n526));
  OAI211_X1 g340(.A(G113), .B(new_n526), .C1(new_n234), .C2(new_n525), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n387), .A2(new_n527), .A3(new_n233), .A4(new_n400), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT81), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n382), .A2(new_n237), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n406), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G122), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n533), .B(KEYINPUT82), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n524), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n535), .ZN(new_n537));
  INV_X1    g351(.A(new_n531), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n391), .B2(new_n396), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n534), .B(new_n523), .C1(new_n539), .C2(new_n530), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n402), .A2(new_n311), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n227), .B2(new_n311), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n190), .A2(G224), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(KEYINPUT7), .B2(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n534), .B(KEYINPUT8), .Z(new_n549));
  AOI21_X1  g363(.A(new_n401), .B1(new_n233), .B2(new_n527), .ZN(new_n550));
  INV_X1    g364(.A(new_n528), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n543), .A2(KEYINPUT7), .A3(new_n547), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n548), .A2(new_n537), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G210), .B1(G237), .B2(G902), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT84), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n559), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AND4_X1   g375(.A1(new_n366), .A2(new_n437), .A3(new_n520), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n310), .A2(new_n359), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT93), .B(G101), .Z(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(G3));
  NOR2_X1   g379(.A1(new_n561), .A2(KEYINPUT94), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT94), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n433), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n432), .A2(new_n436), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n283), .A2(new_n284), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n269), .B2(new_n282), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n359), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n483), .ZN(new_n577));
  INV_X1    g391(.A(new_n366), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n511), .A2(new_n512), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n508), .A2(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT33), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(G478), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n513), .A2(new_n514), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n514), .A2(new_n350), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n577), .A2(new_n578), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  XNOR2_X1  g406(.A(new_n482), .B(KEYINPUT96), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n478), .ZN(new_n594));
  INV_X1    g408(.A(new_n519), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n594), .A2(new_n578), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n576), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT97), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NAND4_X1  g414(.A1(new_n437), .A2(new_n520), .A3(new_n366), .A4(new_n561), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n283), .A2(new_n350), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n344), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT98), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n340), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n355), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n354), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n571), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT37), .B(G110), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  OAI21_X1  g427(.A(new_n362), .B1(new_n364), .B2(G900), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n594), .A2(new_n595), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n310), .A2(new_n570), .A3(new_n616), .A4(new_n609), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT99), .B(G128), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G30));
  NAND2_X1  g433(.A1(new_n304), .A2(new_n194), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n258), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(G472), .B1(new_n621), .B2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n289), .A2(new_n292), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n569), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n614), .B(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT40), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n561), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n483), .B(new_n519), .C1(new_n629), .C2(KEYINPUT40), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n624), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n609), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n433), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT102), .B(G143), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G45));
  NOR3_X1   g453(.A1(new_n577), .A2(new_n588), .A3(new_n615), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n310), .A2(new_n570), .A3(new_n609), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G146), .ZN(G48));
  OR2_X1    g456(.A1(new_n415), .A2(new_n424), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n350), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G469), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n645), .A2(new_n436), .A3(new_n425), .ZN(new_n646));
  INV_X1    g460(.A(new_n568), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n546), .A2(new_n559), .A3(new_n554), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n559), .B1(new_n546), .B2(new_n554), .ZN(new_n649));
  OR3_X1    g463(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT94), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n310), .A3(new_n359), .A4(new_n589), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT41), .B(G113), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G15));
  NAND4_X1  g468(.A1(new_n651), .A2(new_n310), .A3(new_n359), .A4(new_n596), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G116), .ZN(G18));
  NAND3_X1  g470(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT70), .B1(new_n291), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n285), .A2(new_n187), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n636), .B1(new_n660), .B2(new_n309), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n366), .A3(new_n520), .A4(new_n651), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(G472), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n602), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n269), .B1(new_n195), .B2(new_n305), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n284), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n577), .B2(new_n595), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n483), .A2(new_n672), .A3(new_n519), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n651), .A2(new_n670), .A3(new_n674), .A4(new_n366), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  INV_X1    g490(.A(new_n668), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n651), .A2(new_n609), .A3(new_n640), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G125), .ZN(G27));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n285), .B2(new_n288), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n291), .A2(new_n657), .A3(KEYINPUT105), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n309), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n648), .A2(new_n649), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n433), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n569), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n683), .A2(new_n686), .A3(new_n359), .A4(new_n640), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n577), .A2(KEYINPUT42), .A3(new_n588), .A4(new_n615), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n310), .A2(new_n689), .A3(new_n686), .A4(new_n359), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n215), .ZN(G33));
  NAND4_X1  g506(.A1(new_n310), .A2(new_n616), .A3(new_n359), .A4(new_n686), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G134), .ZN(G36));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n636), .B1(new_n603), .B2(new_n571), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n483), .A2(new_n588), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT43), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n685), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n697), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n699), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n428), .A2(new_n429), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT46), .A3(new_n431), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n425), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT46), .B1(new_n708), .B2(new_n431), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n436), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(new_n627), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT108), .B(G137), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT109), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G39));
  OR2_X1    g531(.A1(new_n712), .A2(KEYINPUT47), .ZN(new_n718));
  INV_X1    g532(.A(new_n310), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n712), .A2(KEYINPUT47), .ZN(new_n720));
  INV_X1    g534(.A(new_n685), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(new_n669), .A3(new_n640), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G140), .ZN(G42));
  NOR2_X1   g538(.A1(G952), .A2(G953), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT119), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n360), .A2(G953), .ZN(new_n727));
  INV_X1    g541(.A(new_n646), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n685), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n359), .A2(new_n624), .A3(new_n361), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n588), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n483), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT118), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n632), .A2(new_n728), .A3(new_n433), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n670), .A2(new_n699), .A3(new_n361), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n733), .B(KEYINPUT50), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n736), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(KEYINPUT118), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(KEYINPUT118), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n738), .A2(new_n734), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n729), .A2(new_n699), .A3(new_n361), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n636), .A3(new_n668), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n731), .A2(new_n483), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n746), .B1(new_n730), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n436), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n645), .A2(new_n425), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n718), .A2(new_n720), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n736), .A2(KEYINPUT117), .A3(new_n685), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT117), .B1(new_n736), .B2(new_n685), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n744), .B(new_n748), .C1(new_n751), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT51), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n727), .B(new_n732), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n683), .A2(new_n359), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n745), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT48), .Z(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n661), .B(new_n570), .C1(new_n616), .C2(new_n640), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n609), .A2(new_n615), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n671), .A2(new_n673), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n623), .A3(new_n570), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n766), .A3(new_n678), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n617), .A2(new_n678), .A3(new_n641), .A4(new_n769), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n437), .A2(new_n366), .A3(new_n561), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n595), .A2(new_n483), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n778), .A2(new_n574), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n777), .B1(new_n781), .B2(new_n611), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n684), .A3(new_n578), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n575), .A2(new_n784), .A3(new_n779), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n573), .A2(new_n572), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n290), .A2(new_n287), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(new_n636), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n783), .A2(new_n684), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n366), .A3(new_n520), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n790), .A3(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n782), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT110), .B1(new_n577), .B2(new_n588), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n731), .A2(new_n483), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n575), .A2(new_n797), .A3(new_n784), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n563), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n563), .B2(new_n798), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n662), .B(new_n792), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n686), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n519), .A2(new_n615), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n310), .A2(new_n478), .A3(new_n593), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n677), .A2(new_n640), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n636), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n688), .A2(new_n690), .A3(new_n693), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n652), .A2(new_n655), .A3(new_n675), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n801), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT53), .B1(new_n776), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n800), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n563), .A2(new_n793), .A3(new_n798), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n811), .A2(new_n812), .B1(new_n782), .B2(new_n791), .ZN(new_n813));
  INV_X1    g627(.A(new_n807), .ZN(new_n814));
  INV_X1    g628(.A(new_n808), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n662), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n770), .A2(new_n772), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n806), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n801), .A2(new_n808), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n771), .B(new_n766), .ZN(new_n824));
  INV_X1    g638(.A(new_n806), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n814), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n817), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n809), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT114), .B(KEYINPUT54), .C1(new_n810), .C2(new_n819), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n764), .A2(new_n822), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n738), .A2(new_n651), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n726), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT49), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n669), .B1(new_n750), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n838), .B2(new_n750), .ZN(new_n840));
  INV_X1    g654(.A(new_n433), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(new_n632), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n436), .A3(new_n624), .A4(new_n698), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n843), .ZN(G75));
  NAND2_X1  g658(.A1(new_n360), .A2(G953), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT121), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n350), .B1(new_n827), .B2(new_n830), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n557), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n541), .B(new_n545), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(KEYINPUT55), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(KEYINPUT55), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n853), .B(new_n854), .C1(KEYINPUT120), .C2(new_n850), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(G51));
  AOI211_X1 g672(.A(new_n350), .B(new_n708), .C1(new_n827), .C2(new_n830), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n431), .B(KEYINPUT57), .Z(new_n860));
  AND3_X1   g674(.A1(new_n827), .A2(new_n830), .A3(new_n832), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n832), .B1(new_n827), .B2(new_n830), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n643), .B(KEYINPUT122), .Z(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT123), .B1(new_n865), .B2(new_n847), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n867));
  INV_X1    g681(.A(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n827), .A2(new_n830), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n831), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n833), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n871), .B2(new_n860), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n867), .B(new_n846), .C1(new_n872), .C2(new_n859), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(G54));
  NAND3_X1  g688(.A1(new_n848), .A2(KEYINPUT58), .A3(G475), .ZN(new_n875));
  INV_X1    g689(.A(new_n471), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n847), .B1(new_n877), .B2(new_n878), .ZN(G60));
  NOR2_X1   g693(.A1(new_n582), .A2(new_n583), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n822), .A2(new_n833), .A3(new_n834), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n586), .B(KEYINPUT59), .Z(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n871), .A2(new_n880), .A3(new_n882), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n847), .A3(new_n885), .ZN(G63));
  XNOR2_X1  g700(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n887));
  NAND2_X1  g701(.A1(G217), .A2(G902), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n827), .B2(new_n830), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n847), .B1(new_n890), .B2(new_n607), .ZN(new_n891));
  INV_X1    g705(.A(new_n347), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n890), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G66));
  AOI21_X1  g709(.A(new_n190), .B1(new_n365), .B2(G224), .ZN(new_n896));
  INV_X1    g710(.A(new_n823), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n190), .ZN(new_n898));
  INV_X1    g712(.A(G898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n541), .B1(new_n899), .B2(G953), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n898), .B(new_n900), .ZN(G69));
  XNOR2_X1  g715(.A(new_n257), .B(new_n466), .ZN(new_n902));
  NAND2_X1  g716(.A1(G900), .A2(G953), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n674), .A2(new_n650), .A3(new_n647), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n705), .B1(new_n761), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n713), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n765), .A2(new_n678), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n723), .A3(new_n908), .A4(new_n814), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n902), .B(new_n903), .C1(new_n909), .C2(G953), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n637), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT62), .Z(new_n912));
  NOR3_X1   g726(.A1(new_n719), .A2(new_n669), .A3(new_n802), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n628), .C1(new_n779), .C2(new_n797), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n714), .A3(new_n723), .A4(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n190), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n902), .B(KEYINPUT125), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n910), .B2(KEYINPUT126), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI221_X1 g735(.A(new_n910), .B1(KEYINPUT126), .B2(new_n919), .C1(new_n916), .C2(new_n917), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(G72));
  NAND2_X1  g737(.A1(G472), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT63), .Z(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n915), .B2(new_n897), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n267), .B(KEYINPUT127), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n195), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n909), .B2(new_n897), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n194), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n301), .A2(new_n258), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n925), .B(new_n932), .C1(new_n810), .C2(new_n819), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n846), .A2(new_n929), .A3(new_n931), .A4(new_n933), .ZN(G57));
endmodule


