//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G244), .Z(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  OAI211_X1 g0045(.A(G1), .B(G13), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT68), .A2(G226), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT68), .A2(G226), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT67), .B(G45), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n252), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n244), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n265), .A2(new_n266), .B1(new_n218), .B2(new_n264), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(G222), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n258), .B(new_n260), .C1(new_n272), .C2(new_n246), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT72), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(G200), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n214), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT70), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n205), .A2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G50), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n206), .B1(new_n201), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n244), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n290), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n280), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n287), .B(new_n297), .C1(G50), .C2(new_n283), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT9), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n276), .A2(new_n277), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n273), .A2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G226), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n308), .B(new_n310), .C1(new_n268), .C2(new_n269), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(KEYINPUT82), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n246), .A2(G232), .A3(new_n247), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n256), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G179), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT83), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n311), .A2(KEYINPUT82), .A3(new_n312), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT82), .B1(new_n311), .B2(new_n312), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n325), .A2(new_n326), .A3(new_n246), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n324), .B1(new_n327), .B2(new_n320), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n318), .A2(KEYINPUT83), .A3(new_n321), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n330), .B2(new_n303), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n290), .B1(new_n205), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n285), .A2(new_n332), .B1(new_n284), .B2(new_n290), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n336), .B2(new_n201), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n294), .A2(G159), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n268), .A2(new_n269), .A3(G20), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT79), .B1(new_n341), .B2(KEYINPUT7), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n262), .A2(new_n206), .A3(new_n263), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT79), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n342), .A2(new_n346), .B1(KEYINPUT7), .B2(new_n341), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT16), .B(new_n340), .C1(new_n347), .C2(new_n335), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n279), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT80), .B1(new_n341), .B2(KEYINPUT7), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT80), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n343), .A2(new_n351), .A3(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n263), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT81), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT16), .B1(new_n356), .B2(new_n340), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n333), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n331), .A2(new_n358), .A3(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT84), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n322), .A2(G190), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n330), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n364), .B1(new_n367), .B2(new_n358), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT85), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n246), .B1(new_n313), .B2(new_n314), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n324), .B(new_n320), .C1(new_n370), .C2(new_n316), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT83), .B1(new_n318), .B2(new_n321), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n365), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n333), .ZN(new_n376));
  INV_X1    g0176(.A(new_n279), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n354), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n339), .B1(new_n380), .B2(G68), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n343), .A2(new_n351), .A3(new_n345), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n351), .B1(new_n343), .B2(new_n345), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT81), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n354), .B(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n335), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n383), .B1(new_n389), .B2(new_n339), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n376), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n375), .A2(new_n391), .A3(KEYINPUT84), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n368), .A2(new_n369), .A3(new_n392), .A4(KEYINPUT17), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n368), .A2(KEYINPUT17), .A3(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n375), .A2(new_n391), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT85), .B1(new_n395), .B2(KEYINPUT17), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n363), .B(new_n393), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n264), .A2(G232), .A3(G1698), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n271), .A2(G226), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n317), .ZN(new_n409));
  INV_X1    g0209(.A(new_n256), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(G238), .B2(new_n249), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n398), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n246), .B1(new_n400), .B2(new_n407), .ZN(new_n413));
  INV_X1    g0213(.A(new_n411), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n413), .A2(KEYINPUT13), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(G169), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT14), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(G169), .C1(new_n412), .C2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT75), .B1(new_n413), .B2(new_n414), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n401), .A2(new_n406), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n411), .B(new_n421), .C1(new_n425), .C2(new_n246), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(KEYINPUT13), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G179), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n413), .A2(new_n414), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n398), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n427), .B2(new_n430), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n417), .B(new_n419), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n335), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n288), .B2(new_n295), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n280), .A2(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(KEYINPUT11), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(KEYINPUT11), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT77), .B1(new_n284), .B2(new_n335), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n284), .A2(new_n279), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(G68), .A3(new_n286), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n438), .A2(new_n439), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n434), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G200), .B1(new_n412), .B2(new_n415), .ZN(new_n446));
  INV_X1    g0246(.A(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n415), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n427), .A2(G190), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n449), .A4(G190), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n290), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n458));
  XOR2_X1   g0258(.A(KEYINPUT15), .B(G87), .Z(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n292), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(new_n279), .ZN(new_n462));
  INV_X1    g0262(.A(new_n442), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n286), .A2(G77), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n463), .A2(new_n464), .B1(G77), .B2(new_n283), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n271), .A2(G232), .ZN(new_n467));
  INV_X1    g0267(.A(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G238), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n467), .B1(new_n468), .B2(new_n264), .C1(new_n469), .C2(new_n265), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n317), .ZN(new_n471));
  INV_X1    g0271(.A(new_n217), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n410), .B1(new_n472), .B2(new_n249), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G179), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n466), .B1(new_n475), .B2(KEYINPUT71), .ZN(new_n476));
  AOI21_X1  g0276(.A(G169), .B1(new_n471), .B2(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT71), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(new_n474), .B2(G179), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n462), .A2(new_n465), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n474), .B2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n274), .B2(new_n474), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NOR4_X1   g0284(.A1(new_n306), .A2(new_n397), .A3(new_n456), .A4(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n468), .B1(new_n386), .B2(new_n388), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n468), .A3(KEYINPUT6), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(KEYINPUT6), .B2(new_n488), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT86), .B(G107), .ZN(new_n491));
  XOR2_X1   g0291(.A(new_n490), .B(new_n491), .Z(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n279), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n283), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n205), .A2(G33), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n285), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(G97), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n264), .A2(G244), .A3(new_n307), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT4), .B1(new_n271), .B2(G244), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n317), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n245), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT88), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G41), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(new_n246), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n511), .A3(new_n205), .A4(G45), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n246), .ZN(new_n517));
  INV_X1    g0317(.A(G257), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT89), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT89), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n508), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n366), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G190), .B2(new_n523), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n496), .A2(new_n501), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n303), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G179), .B2(new_n523), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n496), .B2(new_n501), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT90), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n264), .A2(new_n206), .A3(G68), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n292), .A2(new_n488), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(KEYINPUT19), .ZN(new_n534));
  NOR3_X1   g0334(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT19), .B1(new_n404), .B2(new_n405), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(new_n206), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n279), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n460), .A2(new_n284), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n499), .C2(new_n460), .ZN(new_n540));
  INV_X1    g0340(.A(G45), .ZN(new_n541));
  OAI21_X1  g0341(.A(G250), .B1(new_n541), .B2(G1), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n317), .B1(new_n509), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n264), .A2(G244), .A3(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(G238), .B(new_n307), .C1(new_n268), .C2(new_n269), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(G179), .B(new_n543), .C1(new_n547), .C2(new_n317), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n543), .B1(new_n547), .B2(new_n317), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n303), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n366), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n274), .B(new_n543), .C1(new_n547), .C2(new_n317), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n280), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(G87), .A3(new_n283), .A4(new_n498), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n556), .A2(new_n538), .A3(new_n539), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n540), .A2(new_n551), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n530), .A2(new_n531), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n496), .A2(new_n501), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n523), .A2(new_n303), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n523), .A2(G179), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n496), .A2(new_n525), .A3(new_n501), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n558), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n284), .A2(new_n468), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT25), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n499), .B2(new_n468), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n264), .A2(new_n206), .A3(G87), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n468), .A3(G20), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT92), .ZN(new_n578));
  OAI221_X1 g0378(.A(new_n576), .B1(G20), .B2(new_n546), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n578), .B2(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n572), .B1(new_n585), .B2(new_n279), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n264), .A2(G257), .A3(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n264), .A2(G250), .A3(new_n307), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n317), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n516), .A2(new_n246), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G264), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n593), .A3(new_n515), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n303), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G179), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n568), .B1(new_n586), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n498), .A2(G116), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n442), .A2(new_n600), .B1(new_n282), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n503), .B(new_n206), .C1(G33), .C2(new_n488), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT91), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n377), .A2(new_n603), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT20), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n592), .A2(G270), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n264), .A2(G264), .A3(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n264), .A2(G257), .A3(new_n307), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n270), .A2(G303), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n613), .B(new_n515), .C1(new_n617), .C2(new_n246), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G169), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n598), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(G200), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n612), .B(new_n621), .C1(new_n274), .C2(new_n618), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n618), .A2(new_n428), .ZN(new_n623));
  INV_X1    g0423(.A(new_n611), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n604), .B1(new_n624), .B2(new_n609), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(KEYINPUT21), .A3(G169), .A4(new_n618), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n620), .A2(new_n622), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n594), .A2(G200), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n586), .B(new_n629), .C1(new_n274), .C2(new_n594), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n574), .A2(new_n583), .A3(new_n580), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n583), .B1(new_n574), .B2(new_n580), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n279), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n570), .B1(new_n500), .B2(G107), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n596), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT93), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n597), .A2(new_n628), .A3(new_n630), .A4(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n485), .A2(new_n559), .A3(new_n567), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n305), .ZN(new_n640));
  INV_X1    g0440(.A(new_n445), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT95), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n476), .A2(new_n642), .A3(new_n479), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n476), .B2(new_n479), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n455), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n363), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n640), .B1(new_n648), .B2(new_n301), .ZN(new_n649));
  INV_X1    g0449(.A(new_n485), .ZN(new_n650));
  INV_X1    g0450(.A(new_n566), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n620), .A2(new_n626), .A3(new_n627), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n635), .A2(new_n636), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT94), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n630), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n551), .A2(new_n540), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n495), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n490), .B(new_n491), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n660), .A2(new_n206), .B1(new_n218), .B2(new_n295), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(KEYINPUT87), .B2(new_n486), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n377), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n501), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n563), .B(new_n558), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n529), .A2(KEYINPUT26), .A3(new_n558), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n658), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n656), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n649), .B1(new_n650), .B2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n282), .A2(new_n206), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT96), .Z(new_n675));
  INV_X1    g0475(.A(G213), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n673), .B2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n625), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n628), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n620), .A2(new_n626), .A3(new_n627), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n597), .A2(new_n637), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n630), .ZN(new_n687));
  INV_X1    g0487(.A(new_n680), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n586), .A2(new_n688), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n687), .A2(new_n689), .B1(new_n653), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n655), .A2(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(new_n688), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n630), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n535), .A2(new_n601), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n212), .B2(new_n701), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n680), .B1(new_n656), .B2(new_n669), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n597), .A2(new_n683), .A3(new_n637), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n530), .A2(new_n710), .A3(new_n558), .A4(new_n630), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n680), .B1(new_n711), .B2(new_n669), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n708), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n618), .A2(new_n594), .A3(new_n428), .A4(new_n550), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n508), .A2(new_n520), .A3(new_n522), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n317), .A2(new_n590), .B1(new_n592), .B2(G264), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n719), .A2(new_n720), .A3(new_n549), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n719), .B2(new_n549), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n623), .B(new_n716), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT98), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT30), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT30), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n718), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT99), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n559), .A2(new_n567), .A3(new_n638), .A4(new_n688), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n723), .A2(new_n724), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n717), .B1(new_n735), .B2(new_n725), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n680), .B1(new_n736), .B2(KEYINPUT100), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT100), .B(new_n718), .C1(new_n726), .C2(new_n727), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n732), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n730), .A2(new_n731), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n714), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n706), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n281), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n205), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n700), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n685), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G330), .B2(new_n684), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n209), .A2(new_n264), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(KEYINPUT101), .B2(G355), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(KEYINPUT101), .B2(G355), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G116), .B2(new_n209), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n242), .A2(G45), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n209), .A2(new_n270), .ZN(new_n757));
  INV_X1    g0557(.A(new_n255), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(new_n213), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n214), .B1(G20), .B2(new_n303), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n749), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G20), .A3(new_n274), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G329), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n206), .A2(new_n428), .A3(new_n274), .A4(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n270), .B(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n206), .A2(new_n428), .A3(G190), .A4(G200), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT102), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n775), .B1(new_n781), .B2(G311), .ZN(new_n782));
  NAND3_X1  g0582(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(new_n274), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT103), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G326), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n206), .A2(new_n274), .A3(new_n366), .A4(G179), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n206), .B1(new_n768), .B2(G190), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n206), .A2(new_n366), .A3(G179), .A4(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n783), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI22_X1  g0602(.A1(new_n798), .A2(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n782), .A2(new_n790), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT105), .ZN(new_n806));
  INV_X1    g0606(.A(G87), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n264), .B1(new_n792), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n789), .A2(G50), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n781), .A2(G77), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n798), .A2(new_n468), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G68), .B2(new_n800), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n795), .A2(new_n488), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n769), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT104), .B(KEYINPUT32), .Z(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n814), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n816), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(new_n817), .B1(new_n772), .B2(G58), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n811), .A2(new_n813), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n805), .B1(new_n810), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n767), .B1(new_n823), .B2(new_n764), .ZN(new_n824));
  INV_X1    g0624(.A(new_n763), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n684), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n751), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n481), .A2(new_n680), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n645), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n480), .A2(new_n483), .A3(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n707), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n749), .B1(new_n835), .B2(new_n742), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n742), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n749), .ZN(new_n838));
  INV_X1    g0638(.A(new_n764), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n772), .A2(G143), .B1(G150), .B2(new_n800), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n788), .B2(new_n841), .C1(new_n815), .C2(new_n780), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n798), .A2(new_n335), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n270), .B(new_n844), .C1(G132), .C2(new_n770), .ZN(new_n845));
  INV_X1    g0645(.A(new_n795), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n791), .A2(G50), .B1(new_n846), .B2(G58), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G311), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n270), .B1(new_n769), .B2(new_n849), .C1(new_n773), .C2(new_n794), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n781), .B2(G116), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n800), .A2(KEYINPUT106), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n800), .A2(KEYINPUT106), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n789), .A2(G303), .B1(new_n855), .B2(G283), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n798), .A2(new_n807), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n814), .B(new_n857), .C1(G107), .C2(new_n791), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n851), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n839), .B1(new_n848), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n764), .A2(new_n761), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n838), .B(new_n860), .C1(new_n218), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n834), .B2(new_n762), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n837), .A2(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n746), .A2(new_n205), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT100), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n688), .B1(new_n728), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(KEYINPUT31), .A3(new_n738), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n740), .A2(new_n731), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n832), .B1(new_n645), .B2(new_n830), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n444), .A2(new_n680), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n445), .A2(new_n455), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n444), .B(new_n680), .C1(new_n454), .C2(new_n434), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT109), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n555), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT16), .B2(new_n381), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n678), .B1(new_n879), .B2(new_n333), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n397), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n678), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n331), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n333), .B2(new_n879), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n368), .A2(new_n392), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n358), .A2(new_n882), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n359), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n358), .B1(new_n331), .B2(new_n882), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n888), .B1(new_n892), .B2(new_n395), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n375), .A2(new_n391), .A3(KEYINPUT84), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT84), .B1(new_n375), .B2(new_n391), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n359), .A2(new_n887), .A3(new_n888), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT107), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT107), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n885), .A2(new_n889), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n894), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n887), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n902), .A2(KEYINPUT108), .B1(new_n397), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(KEYINPUT107), .A3(new_n898), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n900), .B1(new_n885), .B2(new_n889), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n877), .B1(new_n891), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n881), .B2(new_n890), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(KEYINPUT109), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n875), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n911), .A2(KEYINPUT40), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n485), .A3(new_n869), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n740), .A2(new_n731), .A3(new_n868), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n650), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(G330), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n641), .A2(new_n688), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n902), .A2(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n397), .A2(new_n903), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n909), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n891), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n926), .B(new_n927), .C1(new_n932), .C2(KEYINPUT39), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n363), .A2(new_n882), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n480), .A2(new_n680), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n707), .B2(new_n834), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n872), .A2(new_n873), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n913), .A2(new_n915), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n485), .B1(new_n709), .B2(new_n713), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n649), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n865), .B1(new_n924), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n924), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n492), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n492), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(G116), .A3(new_n215), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n212), .A2(new_n218), .A3(new_n336), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n335), .A2(G50), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n281), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(G367));
  OAI221_X1 g0754(.A(new_n765), .B1(new_n209), .B2(new_n460), .C1(new_n234), .C2(new_n757), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n955), .A2(new_n749), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n657), .A2(new_n688), .A3(new_n557), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n558), .B1(new_n557), .B2(new_n688), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n798), .A2(new_n488), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n270), .B1(new_n769), .B2(new_n961), .C1(new_n773), .C2(new_n793), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(G107), .C2(new_n846), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n799), .B2(new_n780), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n791), .A2(G116), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT46), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n794), .B2(new_n854), .C1(new_n849), .C2(new_n788), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n264), .B1(new_n769), .B2(new_n841), .C1(new_n773), .C2(new_n293), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n781), .B2(G50), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n795), .A2(new_n335), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G77), .B2(new_n797), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n334), .C2(new_n792), .ZN(new_n972));
  INV_X1    g0772(.A(G143), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n788), .A2(new_n973), .B1(new_n854), .B2(new_n815), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n964), .A2(new_n967), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n956), .B1(new_n825), .B2(new_n959), .C1(new_n976), .C2(new_n839), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n560), .A2(new_n680), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n530), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n529), .A2(new_n680), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n696), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n981), .A2(new_n696), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n981), .B2(new_n696), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n685), .A3(new_n690), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(new_n988), .A3(new_n691), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n695), .B1(new_n690), .B2(new_n694), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(new_n685), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n744), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n700), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n748), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n979), .A2(new_n686), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n680), .B1(new_n999), .B2(new_n564), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n981), .A2(new_n695), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n691), .A2(KEYINPUT110), .A3(new_n981), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT110), .B1(new_n691), .B2(new_n981), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1007), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1010));
  OR3_X1    g0810(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1005), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n977), .B1(new_n998), .B2(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(new_n994), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n690), .A2(new_n825), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n231), .A2(new_n758), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1017), .A2(new_n757), .B1(new_n703), .B2(new_n752), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n457), .A2(KEYINPUT50), .A3(new_n288), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT50), .B1(new_n457), .B2(new_n288), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n703), .B(new_n1019), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1018), .A2(new_n1022), .B1(new_n468), .B2(new_n699), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n749), .B1(new_n1023), .B2(new_n766), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n792), .A2(new_n218), .B1(new_n290), .B2(new_n801), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n960), .B(new_n1025), .C1(new_n459), .C2(new_n846), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n789), .A2(G159), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n781), .A2(G68), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n264), .B1(new_n773), .B2(new_n288), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G150), .B2(new_n770), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n264), .B1(new_n770), .B2(G326), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n792), .A2(new_n794), .B1(new_n799), .B2(new_n795), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n781), .A2(G303), .B1(G317), .B2(new_n772), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n849), .B2(new_n854), .C1(new_n774), .C2(new_n788), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1032), .B1(new_n601), .B2(new_n798), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1031), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1024), .B1(new_n1042), .B2(new_n764), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1015), .A2(new_n748), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n744), .A2(new_n1015), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n700), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n744), .A2(new_n1015), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  AND3_X1   g0848(.A1(new_n239), .A2(new_n209), .A3(new_n270), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n765), .B1(new_n488), .B2(new_n209), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n749), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n788), .A2(new_n293), .B1(new_n815), .B2(new_n773), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n792), .A2(new_n335), .B1(new_n218), .B2(new_n795), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n264), .B1(new_n973), .B2(new_n769), .C1(new_n798), .C2(new_n807), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n781), .C2(new_n457), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(new_n288), .C2(new_n854), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n788), .A2(new_n961), .B1(new_n849), .B2(new_n773), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT111), .Z(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n792), .A2(new_n799), .B1(new_n601), .B2(new_n795), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n270), .B1(new_n774), .B2(new_n769), .C1(new_n798), .C2(new_n468), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n781), .C2(G294), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n1063), .C1(new_n793), .C2(new_n854), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1051), .B1(new_n1066), .B2(new_n764), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n981), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n825), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n992), .B2(new_n747), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n990), .A2(new_n991), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n743), .A2(new_n994), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n701), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1045), .A2(new_n992), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  OAI21_X1  g0876(.A(new_n925), .B1(new_n936), .B2(new_n937), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n929), .B1(new_n907), .B2(new_n908), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n902), .A2(KEYINPUT108), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n931), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT39), .B1(new_n1080), .B2(new_n915), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1077), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n935), .B1(new_n712), .B2(new_n834), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n925), .B1(new_n1084), .B2(new_n937), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n932), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT112), .ZN(new_n1089));
  INV_X1    g0889(.A(G330), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n922), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n874), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n927), .B1(new_n932), .B2(KEYINPUT39), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1086), .B1(new_n1095), .B2(new_n1077), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT112), .B1(new_n1096), .B2(new_n1092), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n937), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n741), .A2(new_n1098), .A3(G330), .A4(new_n834), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1083), .A2(new_n1087), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1094), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT113), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n869), .A2(G330), .A3(new_n834), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n937), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1104), .A3(new_n1084), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n741), .A2(G330), .A3(new_n834), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(new_n937), .B1(new_n1091), .B2(new_n874), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1107), .B2(new_n936), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1091), .A2(new_n485), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n942), .A2(new_n1109), .A3(new_n649), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1102), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1101), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1094), .C1(new_n1097), .C2(new_n1100), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n700), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n838), .B1(new_n290), .B2(new_n861), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n844), .B1(G87), .B2(new_n791), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n218), .B2(new_n795), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n780), .A2(new_n488), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n788), .A2(new_n799), .B1(new_n854), .B2(new_n468), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n270), .B1(new_n769), .B2(new_n794), .C1(new_n773), .C2(new_n601), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1124));
  OR3_X1    g0924(.A1(new_n792), .A2(new_n293), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n792), .B2(new_n293), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n772), .A2(G132), .B1(new_n846), .B2(G159), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n264), .B1(new_n1129), .B2(new_n769), .C1(new_n798), .C2(new_n288), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT115), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1128), .B(new_n1131), .C1(G128), .C2(new_n789), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n780), .A2(new_n1133), .B1(new_n841), .B2(new_n854), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT114), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1117), .B1(new_n1136), .B2(new_n839), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1095), .B2(new_n761), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1101), .B2(new_n748), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n1139), .ZN(G378));
  XNOR2_X1  g0940(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n298), .A2(new_n882), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1143));
  OR2_X1    g0943(.A1(new_n306), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n306), .A2(new_n1143), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1141), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1150), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n761), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n772), .A2(G128), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n293), .B2(new_n795), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n800), .A2(G132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n792), .B2(new_n1133), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(new_n781), .C2(G137), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1129), .B2(new_n788), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n797), .A2(G159), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1164));
  AND4_X1   g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n264), .A2(G41), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G50), .B(new_n1166), .C1(new_n244), .C2(new_n245), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n798), .A2(new_n334), .B1(new_n801), .B2(new_n488), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n970), .B(new_n1169), .C1(G77), .C2(new_n791), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1166), .B1(new_n799), .B2(new_n769), .C1(new_n773), .C2(new_n468), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n781), .B2(new_n459), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n601), .C2(new_n788), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT117), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1168), .B1(new_n1174), .B2(KEYINPUT58), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1165), .B(new_n1175), .C1(KEYINPUT58), .C2(new_n1174), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n839), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n838), .B(new_n1177), .C1(new_n288), .C2(new_n861), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1154), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT109), .B1(new_n869), .B2(new_n874), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT40), .B1(new_n932), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n918), .A2(new_n916), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1090), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1183), .A2(new_n941), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n941), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1153), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n933), .B(new_n940), .C1(new_n919), .C2(new_n1090), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n941), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1179), .B1(new_n1191), .B2(new_n747), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(KEYINPUT112), .B(new_n1092), .C1(new_n1083), .C2(new_n1087), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1089), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1108), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1111), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1110), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1190), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n700), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1193), .B1(new_n1201), .B2(new_n1204), .ZN(G375));
  NOR2_X1   g1005(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n997), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n937), .A2(new_n761), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n789), .A2(G132), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n264), .B1(new_n798), .B2(new_n334), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT121), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(KEYINPUT121), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n854), .A2(new_n1133), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n772), .A2(G137), .B1(new_n770), .B2(G128), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G50), .B2(new_n846), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n815), .B2(new_n792), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1217), .B(new_n1221), .C1(G150), .C2(new_n781), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n270), .B1(new_n769), .B2(new_n793), .C1(new_n773), .C2(new_n799), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n846), .A2(new_n459), .B1(new_n797), .B2(G77), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n488), .B2(new_n792), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G107), .C2(new_n781), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n789), .A2(G294), .B1(new_n855), .B2(G116), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1222), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(new_n839), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n838), .B(new_n1229), .C1(new_n335), .C2(new_n861), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1108), .A2(new_n748), .B1(new_n1211), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1209), .A2(new_n1231), .ZN(G381));
  NAND4_X1  g1032(.A1(new_n744), .A2(new_n990), .A3(new_n1015), .A4(new_n991), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n996), .B1(new_n1233), .B2(new_n744), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1011), .B(new_n1012), .C1(new_n1234), .C2(new_n748), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n977), .A3(new_n1075), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n827), .B(new_n1044), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(new_n1209), .A3(new_n1239), .A4(new_n1231), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G378), .A2(G375), .A3(new_n1236), .A4(new_n1240), .ZN(G407));
  NOR2_X1   g1041(.A1(new_n676), .A2(G343), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR3_X1    g1043(.A1(G375), .A2(G378), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G407), .A2(G213), .A3(new_n1244), .ZN(G409));
  NAND2_X1  g1045(.A1(G387), .A2(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT123), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1237), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1247), .B2(new_n1237), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1236), .B(new_n1246), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1237), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1075), .B1(new_n1235), .B2(new_n977), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1255), .A3(KEYINPUT124), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n1250), .C2(new_n1249), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT126), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1193), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1202), .A2(new_n1191), .A3(new_n996), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1116), .B(new_n1139), .C1(new_n1263), .C2(new_n1192), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1243), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1206), .B1(KEYINPUT60), .B2(new_n1208), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1107), .A2(new_n936), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(KEYINPUT60), .A3(new_n1110), .A4(new_n1105), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n700), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1231), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1239), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G384), .B(new_n1231), .C1(new_n1267), .C2(new_n1270), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT122), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1242), .A2(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1272), .A2(new_n1275), .A3(new_n1273), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1276), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1275), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1278), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(new_n1243), .A3(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1261), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1274), .A2(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1265), .A2(new_n1243), .A3(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1242), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1274), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1289), .B1(new_n1296), .B2(new_n1283), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1284), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1260), .B1(new_n1294), .B2(new_n1290), .ZN(new_n1300));
  AND4_X1   g1100(.A1(new_n1289), .A2(new_n1283), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1288), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1304), .B(new_n1288), .C1(new_n1297), .C2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(G405));
  XNOR2_X1  g1106(.A(G375), .B(G378), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1274), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1292), .ZN(G402));
endmodule


