

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n403, n404, n405, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795;

  XNOR2_X1 U380 ( .A(n640), .B(n457), .ZN(n456) );
  AND2_X1 U381 ( .A1(n409), .A2(n407), .ZN(n358) );
  XNOR2_X1 U382 ( .A(n474), .B(KEYINPUT77), .ZN(n692) );
  AND2_X1 U383 ( .A1(n443), .A2(n618), .ZN(n367) );
  NOR2_X1 U384 ( .A1(n752), .A2(G902), .ZN(n518) );
  INV_X1 U385 ( .A(KEYINPUT0), .ZN(n362) );
  XNOR2_X1 U386 ( .A(n359), .B(n565), .ZN(n775) );
  XNOR2_X1 U387 ( .A(n508), .B(G128), .ZN(n563) );
  XNOR2_X1 U388 ( .A(n554), .B(KEYINPUT16), .ZN(n359) );
  XNOR2_X1 U389 ( .A(G101), .B(KEYINPUT66), .ZN(n371) );
  NAND2_X2 U390 ( .A1(n358), .A2(n404), .ZN(n679) );
  XNOR2_X2 U391 ( .A(n543), .B(n365), .ZN(n727) );
  NOR2_X2 U392 ( .A1(n451), .A2(n450), .ZN(n455) );
  XOR2_X2 U393 ( .A(KEYINPUT99), .B(n386), .Z(n590) );
  NAND2_X1 U394 ( .A1(n360), .A2(KEYINPUT47), .ZN(n638) );
  INV_X1 U395 ( .A(n692), .ZN(n360) );
  NAND2_X1 U396 ( .A1(n361), .A2(n462), .ZN(n433) );
  XNOR2_X1 U397 ( .A(n464), .B(n362), .ZN(n361) );
  XNOR2_X2 U398 ( .A(n540), .B(KEYINPUT70), .ZN(n403) );
  NAND2_X2 U399 ( .A1(n382), .A2(n381), .ZN(n540) );
  XNOR2_X1 U400 ( .A(G131), .B(G143), .ZN(n577) );
  INV_X2 U401 ( .A(G953), .ZN(n785) );
  XOR2_X2 U402 ( .A(KEYINPUT40), .B(n611), .Z(n795) );
  XNOR2_X2 U403 ( .A(n384), .B(KEYINPUT0), .ZN(n386) );
  XNOR2_X2 U404 ( .A(n496), .B(KEYINPUT65), .ZN(n657) );
  XOR2_X2 U405 ( .A(KEYINPUT38), .B(n647), .Z(n709) );
  AND2_X1 U406 ( .A1(n650), .A2(n649), .ZN(n783) );
  INV_X1 U407 ( .A(n727), .ZN(n616) );
  OR2_X1 U408 ( .A1(n763), .A2(G902), .ZN(n446) );
  NOR2_X1 U409 ( .A1(n655), .A2(n746), .ZN(n656) );
  AND2_X1 U410 ( .A1(n485), .A2(n484), .ZN(n481) );
  AND2_X1 U411 ( .A1(n491), .A2(n490), .ZN(n489) );
  XNOR2_X1 U412 ( .A(n420), .B(n418), .ZN(n763) );
  INV_X1 U413 ( .A(G143), .ZN(n508) );
  NOR2_X2 U414 ( .A1(n657), .A2(n656), .ZN(n761) );
  XNOR2_X1 U415 ( .A(n475), .B(n370), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n617), .B(n519), .ZN(n644) );
  XNOR2_X1 U417 ( .A(KEYINPUT33), .B(KEYINPUT90), .ZN(n544) );
  INV_X1 U418 ( .A(KEYINPUT78), .ZN(n394) );
  NOR2_X1 U419 ( .A1(G953), .A2(G237), .ZN(n573) );
  XNOR2_X1 U420 ( .A(n563), .B(n509), .ZN(n550) );
  INV_X1 U421 ( .A(KEYINPUT4), .ZN(n509) );
  NOR2_X1 U422 ( .A1(n672), .A2(G902), .ZN(n543) );
  XNOR2_X1 U423 ( .A(n440), .B(n439), .ZN(n642) );
  INV_X1 U424 ( .A(KEYINPUT39), .ZN(n439) );
  NOR2_X1 U425 ( .A1(n635), .A2(n610), .ZN(n440) );
  AND2_X1 U426 ( .A1(n714), .A2(n473), .ZN(n472) );
  INV_X1 U427 ( .A(KEYINPUT47), .ZN(n473) );
  INV_X1 U428 ( .A(KEYINPUT79), .ZN(n457) );
  AND2_X1 U429 ( .A1(n480), .A2(n413), .ZN(n393) );
  AND2_X1 U430 ( .A1(n480), .A2(n588), .ZN(n423) );
  AND2_X1 U431 ( .A1(n481), .A2(n413), .ZN(n389) );
  INV_X1 U432 ( .A(KEYINPUT67), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n460), .B(n459), .ZN(n562) );
  XNOR2_X1 U434 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n459) );
  XNOR2_X1 U435 ( .A(n461), .B(KEYINPUT68), .ZN(n460) );
  NAND2_X1 U436 ( .A1(n785), .A2(G234), .ZN(n461) );
  XNOR2_X1 U437 ( .A(n479), .B(G122), .ZN(n565) );
  XNOR2_X1 U438 ( .A(G116), .B(G107), .ZN(n479) );
  XNOR2_X1 U439 ( .A(n553), .B(n550), .ZN(n400) );
  XNOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT95), .ZN(n551) );
  XOR2_X1 U441 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n552) );
  NOR2_X1 U442 ( .A1(n561), .A2(n494), .ZN(n490) );
  AND2_X1 U443 ( .A1(n619), .A2(n495), .ZN(n494) );
  INV_X1 U444 ( .A(KEYINPUT1), .ZN(n519) );
  XNOR2_X1 U445 ( .A(n781), .B(n471), .ZN(n672) );
  XNOR2_X1 U446 ( .A(n441), .B(n542), .ZN(n471) );
  XNOR2_X1 U447 ( .A(n536), .B(n541), .ZN(n441) );
  XOR2_X1 U448 ( .A(G110), .B(G137), .Z(n530) );
  XNOR2_X1 U449 ( .A(G119), .B(G128), .ZN(n529) );
  XNOR2_X1 U450 ( .A(n527), .B(n422), .ZN(n421) );
  XNOR2_X1 U451 ( .A(n528), .B(KEYINPUT23), .ZN(n422) );
  XNOR2_X1 U452 ( .A(KEYINPUT10), .B(G140), .ZN(n419) );
  XNOR2_X1 U453 ( .A(G134), .B(KEYINPUT108), .ZN(n438) );
  XNOR2_X1 U454 ( .A(n535), .B(n470), .ZN(n469) );
  XNOR2_X1 U455 ( .A(n511), .B(G107), .ZN(n470) );
  INV_X1 U456 ( .A(KEYINPUT32), .ZN(n486) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n607) );
  INV_X1 U458 ( .A(KEYINPUT30), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n445), .B(n444), .ZN(n443) );
  INV_X1 U460 ( .A(KEYINPUT28), .ZN(n444) );
  OR2_X1 U461 ( .A1(n619), .A2(n495), .ZN(n493) );
  XNOR2_X1 U462 ( .A(n433), .B(KEYINPUT22), .ZN(n585) );
  AND2_X1 U463 ( .A1(n711), .A2(n724), .ZN(n462) );
  NOR2_X1 U464 ( .A1(n412), .A2(n411), .ZN(n410) );
  NOR2_X1 U465 ( .A1(n722), .A2(KEYINPUT87), .ZN(n408) );
  INV_X1 U466 ( .A(KEYINPUT87), .ZN(n411) );
  XOR2_X1 U467 ( .A(KEYINPUT93), .B(n664), .Z(n765) );
  NAND2_X1 U468 ( .A1(n456), .A2(KEYINPUT72), .ZN(n447) );
  AND2_X1 U469 ( .A1(n449), .A2(n702), .ZN(n448) );
  AND2_X1 U470 ( .A1(n452), .A2(n453), .ZN(n451) );
  OR2_X1 U471 ( .A1(G237), .A2(G902), .ZN(n547) );
  XOR2_X1 U472 ( .A(KEYINPUT103), .B(KEYINPUT20), .Z(n521) );
  XNOR2_X1 U473 ( .A(G116), .B(KEYINPUT74), .ZN(n537) );
  XOR2_X1 U474 ( .A(KEYINPUT5), .B(KEYINPUT105), .Z(n538) );
  NAND2_X1 U475 ( .A1(n454), .A2(n455), .ZN(n436) );
  XNOR2_X1 U476 ( .A(n458), .B(n624), .ZN(n454) );
  NAND2_X1 U477 ( .A1(n447), .A2(n448), .ZN(n450) );
  INV_X1 U478 ( .A(KEYINPUT48), .ZN(n435) );
  XNOR2_X1 U479 ( .A(n535), .B(G131), .ZN(n781) );
  XNOR2_X1 U480 ( .A(n475), .B(n370), .ZN(n770) );
  XNOR2_X1 U481 ( .A(KEYINPUT80), .B(KEYINPUT101), .ZN(n525) );
  XNOR2_X1 U482 ( .A(G113), .B(G104), .ZN(n570) );
  XOR2_X1 U483 ( .A(KEYINPUT12), .B(KEYINPUT106), .Z(n575) );
  XNOR2_X1 U484 ( .A(G146), .B(G131), .ZN(n511) );
  XNOR2_X1 U485 ( .A(n516), .B(n503), .ZN(n502) );
  INV_X1 U486 ( .A(G140), .ZN(n503) );
  XNOR2_X1 U487 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U488 ( .A(KEYINPUT76), .ZN(n514) );
  XNOR2_X1 U489 ( .A(n550), .B(n510), .ZN(n535) );
  XNOR2_X1 U490 ( .A(G137), .B(G134), .ZN(n510) );
  NAND2_X1 U491 ( .A1(G234), .A2(G237), .ZN(n556) );
  XNOR2_X1 U492 ( .A(KEYINPUT111), .B(n620), .ZN(n715) );
  XNOR2_X1 U493 ( .A(n727), .B(KEYINPUT6), .ZN(n628) );
  XNOR2_X1 U494 ( .A(n513), .B(G110), .ZN(n773) );
  XNOR2_X1 U495 ( .A(G104), .B(KEYINPUT94), .ZN(n513) );
  XNOR2_X1 U496 ( .A(n400), .B(n399), .ZN(n398) );
  XNOR2_X1 U497 ( .A(n549), .B(n366), .ZN(n399) );
  XNOR2_X1 U498 ( .A(n507), .B(n782), .ZN(n418) );
  XNOR2_X1 U499 ( .A(n531), .B(n421), .ZN(n420) );
  XNOR2_X1 U500 ( .A(n567), .B(n437), .ZN(n759) );
  XNOR2_X1 U501 ( .A(n568), .B(n566), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n563), .B(n438), .ZN(n564) );
  XNOR2_X1 U503 ( .A(n666), .B(n665), .ZN(n667) );
  INV_X1 U504 ( .A(n634), .ZN(n465) );
  NAND2_X1 U505 ( .A1(n722), .A2(n486), .ZN(n484) );
  NAND2_X1 U506 ( .A1(n483), .A2(n482), .ZN(n480) );
  NOR2_X1 U507 ( .A1(n722), .A2(n486), .ZN(n482) );
  NOR2_X1 U508 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U509 ( .A1(n367), .A2(n364), .ZN(n474) );
  NOR2_X1 U510 ( .A1(n597), .A2(n596), .ZN(n686) );
  NAND2_X1 U511 ( .A1(n722), .A2(n415), .ZN(n414) );
  NOR2_X1 U512 ( .A1(n408), .A2(n586), .ZN(n407) );
  NAND2_X1 U513 ( .A1(n405), .A2(n411), .ZN(n404) );
  XNOR2_X1 U514 ( .A(n673), .B(KEYINPUT62), .ZN(n674) );
  XNOR2_X1 U515 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U516 ( .A(n754), .B(n753), .ZN(n755) );
  INV_X1 U517 ( .A(KEYINPUT56), .ZN(n504) );
  AND2_X1 U518 ( .A1(n368), .A2(n492), .ZN(n364) );
  XOR2_X1 U519 ( .A(G472), .B(KEYINPUT71), .Z(n365) );
  AND2_X1 U520 ( .A1(G224), .A2(n785), .ZN(n366) );
  INV_X1 U521 ( .A(n413), .ZN(n685) );
  AND2_X1 U522 ( .A1(n491), .A2(n488), .ZN(n368) );
  AND2_X1 U523 ( .A1(n481), .A2(n480), .ZN(n369) );
  XOR2_X1 U524 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n370) );
  INV_X1 U525 ( .A(n588), .ZN(n487) );
  INV_X1 U526 ( .A(KEYINPUT82), .ZN(n432) );
  XNOR2_X1 U527 ( .A(G101), .B(KEYINPUT66), .ZN(n512) );
  XNOR2_X1 U528 ( .A(n395), .B(n394), .ZN(n639) );
  NAND2_X1 U529 ( .A1(n690), .A2(n434), .ZN(n395) );
  NAND2_X1 U530 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U531 ( .A(n372), .B(KEYINPUT73), .ZN(n641) );
  NAND2_X1 U532 ( .A1(n692), .A2(n472), .ZN(n372) );
  NOR2_X1 U533 ( .A1(n616), .A2(n725), .ZN(n415) );
  NAND2_X1 U534 ( .A1(n725), .A2(n724), .ZN(n721) );
  NOR2_X1 U535 ( .A1(n725), .A2(n615), .ZN(n625) );
  NAND2_X1 U536 ( .A1(n661), .A2(n651), .ZN(n373) );
  NAND2_X1 U537 ( .A1(n775), .A2(n424), .ZN(n376) );
  NAND2_X1 U538 ( .A1(n374), .A2(n375), .ZN(n377) );
  NAND2_X1 U539 ( .A1(n376), .A2(n377), .ZN(n401) );
  INV_X1 U540 ( .A(n775), .ZN(n374) );
  INV_X1 U541 ( .A(n424), .ZN(n375) );
  BUF_X1 U542 ( .A(n661), .Z(n378) );
  NAND2_X1 U543 ( .A1(n371), .A2(KEYINPUT67), .ZN(n381) );
  NAND2_X1 U544 ( .A1(n379), .A2(n380), .ZN(n382) );
  INV_X1 U545 ( .A(n512), .ZN(n379) );
  NAND2_X1 U546 ( .A1(n661), .A2(n651), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n442), .B(n555), .ZN(n383) );
  XNOR2_X1 U548 ( .A(n373), .B(n555), .ZN(n629) );
  OR2_X1 U549 ( .A1(n585), .A2(n414), .ZN(n413) );
  XNOR2_X2 U550 ( .A(n622), .B(KEYINPUT42), .ZN(n794) );
  INV_X1 U551 ( .A(n383), .ZN(n647) );
  XNOR2_X1 U552 ( .A(n436), .B(n435), .ZN(n650) );
  NAND2_X1 U553 ( .A1(n416), .A2(n628), .ZN(n545) );
  XNOR2_X1 U554 ( .A(n592), .B(KEYINPUT110), .ZN(n416) );
  NAND2_X1 U555 ( .A1(n492), .A2(n489), .ZN(n384) );
  NAND2_X1 U556 ( .A1(n489), .A2(n492), .ZN(n464) );
  XNOR2_X2 U557 ( .A(KEYINPUT41), .B(n621), .ZN(n737) );
  NOR2_X1 U558 ( .A1(n657), .A2(n656), .ZN(n385) );
  INV_X1 U559 ( .A(n647), .ZN(n387) );
  BUF_X1 U560 ( .A(n363), .Z(n388) );
  OR2_X2 U561 ( .A1(n792), .A2(KEYINPUT44), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n517), .B(n469), .ZN(n752) );
  NAND2_X1 U563 ( .A1(n423), .A2(n389), .ZN(n390) );
  NAND2_X1 U564 ( .A1(n391), .A2(n390), .ZN(n589) );
  NAND2_X1 U565 ( .A1(n392), .A2(n487), .ZN(n391) );
  NAND2_X1 U566 ( .A1(n393), .A2(n481), .ZN(n392) );
  NAND2_X1 U567 ( .A1(n679), .A2(n601), .ZN(n498) );
  NAND2_X1 U568 ( .A1(n608), .A2(n609), .ZN(n635) );
  NOR2_X1 U569 ( .A1(n727), .A2(n619), .ZN(n397) );
  XNOR2_X2 U570 ( .A(n446), .B(n532), .ZN(n586) );
  XNOR2_X2 U571 ( .A(n401), .B(n398), .ZN(n661) );
  XNOR2_X2 U572 ( .A(n403), .B(n773), .ZN(n424) );
  INV_X1 U573 ( .A(n600), .ZN(n405) );
  NAND2_X1 U574 ( .A1(n600), .A2(n410), .ZN(n409) );
  INV_X1 U575 ( .A(n722), .ZN(n412) );
  AND2_X2 U576 ( .A1(n417), .A2(n644), .ZN(n592) );
  INV_X1 U577 ( .A(n721), .ZN(n417) );
  XNOR2_X1 U578 ( .A(n548), .B(n419), .ZN(n782) );
  XNOR2_X1 U579 ( .A(n369), .B(G119), .ZN(G21) );
  XNOR2_X1 U580 ( .A(n424), .B(n502), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n770), .A2(KEYINPUT82), .ZN(n428) );
  NAND2_X1 U582 ( .A1(n425), .A2(n783), .ZN(n497) );
  NOR2_X1 U583 ( .A1(n426), .A2(n429), .ZN(n425) );
  NAND2_X1 U584 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U585 ( .A1(n651), .A2(KEYINPUT82), .ZN(n427) );
  NOR2_X1 U586 ( .A1(n363), .A2(n430), .ZN(n429) );
  NAND2_X1 U587 ( .A1(n431), .A2(n432), .ZN(n430) );
  INV_X1 U588 ( .A(n651), .ZN(n431) );
  XNOR2_X2 U589 ( .A(n583), .B(KEYINPUT35), .ZN(n792) );
  NAND2_X1 U590 ( .A1(n633), .A2(KEYINPUT47), .ZN(n434) );
  OR2_X2 U591 ( .A1(n383), .A2(n493), .ZN(n492) );
  INV_X1 U592 ( .A(n590), .ZN(n501) );
  NAND2_X1 U593 ( .A1(n625), .A2(n616), .ZN(n445) );
  NAND2_X1 U594 ( .A1(n641), .A2(KEYINPUT72), .ZN(n449) );
  INV_X1 U595 ( .A(n456), .ZN(n453) );
  NOR2_X1 U596 ( .A1(n641), .A2(KEYINPUT72), .ZN(n452) );
  NAND2_X1 U597 ( .A1(n795), .A2(n794), .ZN(n458) );
  AND2_X2 U598 ( .A1(n466), .A2(n465), .ZN(n583) );
  XNOR2_X1 U599 ( .A(n468), .B(n467), .ZN(n466) );
  INV_X1 U600 ( .A(KEYINPUT34), .ZN(n467) );
  NAND2_X1 U601 ( .A1(n706), .A2(n501), .ZN(n468) );
  XNOR2_X2 U602 ( .A(n545), .B(n544), .ZN(n706) );
  INV_X1 U603 ( .A(n644), .ZN(n722) );
  INV_X2 U604 ( .A(n586), .ZN(n725) );
  XNOR2_X1 U605 ( .A(n498), .B(KEYINPUT109), .ZN(n476) );
  NAND2_X1 U606 ( .A1(n647), .A2(n636), .ZN(n690) );
  NOR2_X1 U607 ( .A1(n612), .A2(n607), .ZN(n608) );
  NAND2_X1 U608 ( .A1(n497), .A2(n653), .ZN(n496) );
  NAND2_X1 U609 ( .A1(n477), .A2(n476), .ZN(n475) );
  NAND2_X1 U610 ( .A1(n499), .A2(n500), .ZN(n477) );
  XNOR2_X2 U611 ( .A(n478), .B(G119), .ZN(n554) );
  XNOR2_X2 U612 ( .A(G113), .B(KEYINPUT3), .ZN(n478) );
  INV_X1 U613 ( .A(n587), .ZN(n483) );
  NAND2_X1 U614 ( .A1(n587), .A2(n486), .ZN(n485) );
  INV_X1 U615 ( .A(n494), .ZN(n488) );
  NAND2_X1 U616 ( .A1(n629), .A2(n495), .ZN(n491) );
  INV_X1 U617 ( .A(KEYINPUT19), .ZN(n495) );
  NAND2_X1 U618 ( .A1(n589), .A2(n792), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n505), .B(n504), .ZN(G51) );
  NAND2_X1 U620 ( .A1(n506), .A2(n676), .ZN(n505) );
  XNOR2_X1 U621 ( .A(n663), .B(n662), .ZN(n506) );
  XOR2_X1 U622 ( .A(n530), .B(n529), .Z(n507) );
  XOR2_X1 U623 ( .A(G146), .B(G125), .Z(n548) );
  INV_X1 U624 ( .A(n548), .ZN(n549) );
  XNOR2_X1 U625 ( .A(n554), .B(G146), .ZN(n536) );
  INV_X1 U626 ( .A(n703), .ZN(n648) );
  INV_X1 U627 ( .A(KEYINPUT100), .ZN(n528) );
  NOR2_X1 U628 ( .A1(n648), .A2(n705), .ZN(n649) );
  XNOR2_X1 U629 ( .A(n675), .B(n674), .ZN(n677) );
  XNOR2_X1 U630 ( .A(n668), .B(n667), .ZN(n669) );
  INV_X1 U631 ( .A(KEYINPUT60), .ZN(n670) );
  NAND2_X1 U632 ( .A1(G227), .A2(n785), .ZN(n515) );
  XNOR2_X2 U633 ( .A(n518), .B(G469), .ZN(n617) );
  XOR2_X1 U634 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n523) );
  XNOR2_X2 U635 ( .A(G902), .B(KEYINPUT15), .ZN(n651) );
  NAND2_X1 U636 ( .A1(G234), .A2(n651), .ZN(n520) );
  XNOR2_X1 U637 ( .A(n521), .B(n520), .ZN(n533) );
  NAND2_X1 U638 ( .A1(G217), .A2(n533), .ZN(n522) );
  XNOR2_X1 U639 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U640 ( .A(KEYINPUT104), .B(n524), .ZN(n532) );
  XOR2_X1 U641 ( .A(KEYINPUT102), .B(KEYINPUT24), .Z(n526) );
  XNOR2_X1 U642 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U643 ( .A1(n562), .A2(G221), .ZN(n531) );
  NAND2_X1 U644 ( .A1(G221), .A2(n533), .ZN(n534) );
  XOR2_X1 U645 ( .A(n534), .B(KEYINPUT21), .Z(n724) );
  XNOR2_X1 U646 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U647 ( .A(n540), .B(n539), .Z(n542) );
  NAND2_X1 U648 ( .A1(n573), .A2(G210), .ZN(n541) );
  NAND2_X1 U649 ( .A1(n547), .A2(G214), .ZN(n546) );
  XOR2_X1 U650 ( .A(n546), .B(KEYINPUT96), .Z(n619) );
  NAND2_X1 U651 ( .A1(G210), .A2(n547), .ZN(n555) );
  XNOR2_X1 U652 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U653 ( .A(G898), .B(KEYINPUT97), .ZN(n768) );
  NAND2_X1 U654 ( .A1(G953), .A2(n768), .ZN(n776) );
  XOR2_X1 U655 ( .A(n556), .B(KEYINPUT14), .Z(n742) );
  INV_X1 U656 ( .A(n742), .ZN(n605) );
  NAND2_X1 U657 ( .A1(G902), .A2(n605), .ZN(n557) );
  NOR2_X1 U658 ( .A1(n776), .A2(n557), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n558), .B(KEYINPUT98), .ZN(n560) );
  NAND2_X1 U660 ( .A1(G952), .A2(n785), .ZN(n603) );
  NOR2_X1 U661 ( .A1(n603), .A2(n742), .ZN(n559) );
  NOR2_X1 U662 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U663 ( .A1(G217), .A2(n562), .ZN(n568) );
  XOR2_X1 U664 ( .A(n564), .B(KEYINPUT9), .Z(n567) );
  XNOR2_X1 U665 ( .A(n565), .B(KEYINPUT7), .ZN(n566) );
  NOR2_X1 U666 ( .A1(G902), .A2(n759), .ZN(n569) );
  XOR2_X1 U667 ( .A(G478), .B(n569), .Z(n595) );
  XNOR2_X1 U668 ( .A(KEYINPUT13), .B(G475), .ZN(n582) );
  XOR2_X1 U669 ( .A(KEYINPUT107), .B(G122), .Z(n571) );
  XNOR2_X1 U670 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n782), .B(n572), .ZN(n580) );
  NAND2_X1 U672 ( .A1(G214), .A2(n573), .ZN(n574) );
  XNOR2_X1 U673 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U674 ( .A(n576), .B(KEYINPUT11), .Z(n578) );
  XNOR2_X1 U675 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U676 ( .A(n580), .B(n579), .ZN(n666) );
  NOR2_X1 U677 ( .A1(G902), .A2(n666), .ZN(n581) );
  XNOR2_X1 U678 ( .A(n582), .B(n581), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n595), .A2(n597), .ZN(n634) );
  INV_X1 U680 ( .A(KEYINPUT44), .ZN(n584) );
  NAND2_X1 U681 ( .A1(n584), .A2(KEYINPUT88), .ZN(n588) );
  NOR2_X1 U682 ( .A1(n595), .A2(n597), .ZN(n711) );
  INV_X1 U683 ( .A(n724), .ZN(n613) );
  NOR2_X2 U684 ( .A1(n585), .A2(n628), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n599), .A2(n586), .ZN(n587) );
  NOR2_X1 U686 ( .A1(n721), .A2(n617), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n616), .A2(n590), .ZN(n591) );
  NAND2_X1 U688 ( .A1(n609), .A2(n591), .ZN(n681) );
  NAND2_X1 U689 ( .A1(n616), .A2(n592), .ZN(n733) );
  NOR2_X1 U690 ( .A1(n733), .A2(n386), .ZN(n594) );
  XNOR2_X1 U691 ( .A(n594), .B(KEYINPUT31), .ZN(n697) );
  NAND2_X1 U692 ( .A1(n681), .A2(n697), .ZN(n598) );
  INV_X1 U693 ( .A(n595), .ZN(n596) );
  INV_X1 U694 ( .A(n686), .ZN(n698) );
  NAND2_X1 U695 ( .A1(n597), .A2(n596), .ZN(n694) );
  NAND2_X1 U696 ( .A1(n698), .A2(n694), .ZN(n714) );
  NAND2_X1 U697 ( .A1(n598), .A2(n714), .ZN(n601) );
  XNOR2_X1 U698 ( .A(n599), .B(KEYINPUT86), .ZN(n600) );
  INV_X1 U699 ( .A(n709), .ZN(n610) );
  NOR2_X1 U700 ( .A1(G900), .A2(n785), .ZN(n602) );
  NAND2_X1 U701 ( .A1(n602), .A2(G902), .ZN(n604) );
  NAND2_X1 U702 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U703 ( .A1(n606), .A2(n605), .ZN(n612) );
  INV_X1 U704 ( .A(n694), .ZN(n691) );
  AND2_X1 U705 ( .A1(n642), .A2(n691), .ZN(n611) );
  NOR2_X1 U706 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U707 ( .A(n614), .B(KEYINPUT69), .ZN(n615) );
  INV_X1 U708 ( .A(n617), .ZN(n618) );
  INV_X1 U709 ( .A(n619), .ZN(n708) );
  NAND2_X1 U710 ( .A1(n709), .A2(n708), .ZN(n620) );
  NAND2_X1 U711 ( .A1(n715), .A2(n711), .ZN(n621) );
  NAND2_X1 U712 ( .A1(n367), .A2(n737), .ZN(n622) );
  XNOR2_X1 U713 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n623) );
  XNOR2_X1 U714 ( .A(n623), .B(KEYINPUT64), .ZN(n624) );
  XOR2_X1 U715 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n631) );
  NAND2_X1 U716 ( .A1(n708), .A2(n625), .ZN(n626) );
  NOR2_X1 U717 ( .A1(n694), .A2(n626), .ZN(n627) );
  NAND2_X1 U718 ( .A1(n628), .A2(n627), .ZN(n643) );
  OR2_X1 U719 ( .A1(n643), .A2(n387), .ZN(n630) );
  XNOR2_X1 U720 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U721 ( .A1(n632), .A2(n412), .ZN(n702) );
  INV_X1 U722 ( .A(n714), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n686), .A2(n642), .ZN(n703) );
  NOR2_X1 U724 ( .A1(n412), .A2(n643), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(KEYINPUT43), .ZN(n646) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n705) );
  XNOR2_X1 U727 ( .A(n651), .B(KEYINPUT83), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  INV_X1 U729 ( .A(KEYINPUT2), .ZN(n655) );
  INV_X1 U730 ( .A(n388), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n783), .A2(n654), .ZN(n746) );
  NAND2_X1 U732 ( .A1(n761), .A2(G210), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT89), .B(KEYINPUT55), .Z(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U736 ( .A(n378), .B(n660), .Z(n662) );
  NOR2_X1 U737 ( .A1(G952), .A2(n785), .ZN(n664) );
  INV_X1 U738 ( .A(n765), .ZN(n676) );
  NAND2_X1 U739 ( .A1(n761), .A2(G475), .ZN(n668) );
  XOR2_X1 U740 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n665) );
  NAND2_X1 U741 ( .A1(n669), .A2(n676), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n761), .A2(G472), .ZN(n675) );
  XOR2_X1 U744 ( .A(n672), .B(KEYINPUT92), .Z(n673) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U747 ( .A(n679), .B(G101), .ZN(G3) );
  NOR2_X1 U748 ( .A1(n694), .A2(n681), .ZN(n680) );
  XOR2_X1 U749 ( .A(G104), .B(n680), .Z(G6) );
  NOR2_X1 U750 ( .A1(n698), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U753 ( .A(G107), .B(n684), .ZN(G9) );
  XOR2_X1 U754 ( .A(G110), .B(n685), .Z(G12) );
  XOR2_X1 U755 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U756 ( .A1(n692), .A2(n686), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U758 ( .A(G128), .B(n689), .Z(G30) );
  XNOR2_X1 U759 ( .A(G143), .B(n690), .ZN(G45) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n693), .B(G146), .ZN(G48) );
  NOR2_X1 U762 ( .A1(n694), .A2(n697), .ZN(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(n695), .Z(n696) );
  XNOR2_X1 U764 ( .A(G113), .B(n696), .ZN(G15) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U766 ( .A(G116), .B(KEYINPUT115), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n700), .B(n699), .ZN(G18) );
  XOR2_X1 U768 ( .A(G125), .B(KEYINPUT37), .Z(n701) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(KEYINPUT116), .ZN(n704) );
  XNOR2_X1 U771 ( .A(n704), .B(n703), .ZN(G36) );
  XOR2_X1 U772 ( .A(G140), .B(n705), .Z(G42) );
  BUF_X1 U773 ( .A(n706), .Z(n719) );
  NAND2_X1 U774 ( .A1(n737), .A2(n719), .ZN(n707) );
  XNOR2_X1 U775 ( .A(n707), .B(KEYINPUT122), .ZN(n745) );
  NOR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U777 ( .A(KEYINPUT119), .B(n710), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT120), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U783 ( .A(KEYINPUT121), .B(n720), .Z(n739) );
  NAND2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U785 ( .A(KEYINPUT50), .B(n723), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U787 ( .A(n726), .B(KEYINPUT49), .ZN(n728) );
  NAND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U789 ( .A(KEYINPUT117), .B(n729), .ZN(n730) );
  NAND2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U791 ( .A(n732), .B(KEYINPUT118), .ZN(n734) );
  NAND2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U793 ( .A(KEYINPUT51), .B(n735), .Z(n736) );
  NAND2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U796 ( .A(KEYINPUT52), .B(n740), .Z(n741) );
  NOR2_X1 U797 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n743), .A2(G952), .ZN(n744) );
  NAND2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n748) );
  XNOR2_X1 U800 ( .A(KEYINPUT2), .B(n746), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(KEYINPUT123), .ZN(n750) );
  NOR2_X1 U803 ( .A1(G953), .A2(n750), .ZN(n751) );
  XNOR2_X1 U804 ( .A(KEYINPUT53), .B(n751), .ZN(G75) );
  NAND2_X1 U805 ( .A1(n385), .A2(G469), .ZN(n756) );
  BUF_X1 U806 ( .A(n752), .Z(n754) );
  XOR2_X1 U807 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n753) );
  NOR2_X1 U808 ( .A1(n765), .A2(n757), .ZN(G54) );
  NAND2_X1 U809 ( .A1(G478), .A2(n385), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n765), .A2(n760), .ZN(G63) );
  NAND2_X1 U812 ( .A1(G217), .A2(n385), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U814 ( .A1(n765), .A2(n764), .ZN(G66) );
  XOR2_X1 U815 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n767) );
  NAND2_X1 U816 ( .A1(G224), .A2(G953), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n767), .B(n766), .ZN(n769) );
  NOR2_X1 U818 ( .A1(n769), .A2(n768), .ZN(n772) );
  NOR2_X1 U819 ( .A1(G953), .A2(n388), .ZN(n771) );
  NOR2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n779) );
  XOR2_X1 U821 ( .A(n773), .B(G101), .Z(n774) );
  XNOR2_X1 U822 ( .A(n775), .B(n774), .ZN(n777) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U824 ( .A(n779), .B(n778), .Z(n780) );
  XNOR2_X1 U825 ( .A(KEYINPUT127), .B(n780), .ZN(G69) );
  XOR2_X1 U826 ( .A(n782), .B(n781), .Z(n787) );
  INV_X1 U827 ( .A(n787), .ZN(n784) );
  XOR2_X1 U828 ( .A(n784), .B(n783), .Z(n786) );
  NAND2_X1 U829 ( .A1(n786), .A2(n785), .ZN(n791) );
  XOR2_X1 U830 ( .A(G227), .B(n787), .Z(n788) );
  NAND2_X1 U831 ( .A1(n788), .A2(G900), .ZN(n789) );
  NAND2_X1 U832 ( .A1(n789), .A2(G953), .ZN(n790) );
  NAND2_X1 U833 ( .A1(n791), .A2(n790), .ZN(G72) );
  INV_X1 U834 ( .A(n792), .ZN(n793) );
  XOR2_X1 U835 ( .A(G122), .B(n793), .Z(G24) );
  XNOR2_X1 U836 ( .A(G137), .B(n794), .ZN(G39) );
  XNOR2_X1 U837 ( .A(G131), .B(n795), .ZN(G33) );
endmodule

