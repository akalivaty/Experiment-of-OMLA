//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n213), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n221), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT67), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT70), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n209), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT72), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n217), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n208), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G50), .B2(new_n264), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n275), .A2(G223), .B1(G77), .B2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(G222), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G1), .A2(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G41), .A2(G45), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT71), .B1(new_n290), .B2(G1), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n208), .C1(G41), .C2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n285), .B2(new_n286), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n208), .A2(new_n301), .B1(new_n285), .B2(new_n286), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(G226), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n289), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n270), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n289), .A2(new_n307), .A3(new_n303), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(new_n270), .B(KEYINPUT9), .Z(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G200), .B2(new_n304), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(G200), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n311), .A3(new_n314), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n310), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n257), .A2(new_n253), .B1(new_n209), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n255), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n261), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n327), .B(KEYINPUT73), .Z(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n208), .B2(G20), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n266), .A2(new_n329), .B1(new_n323), .B2(new_n265), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n275), .A2(G238), .B1(G107), .B2(new_n273), .ZN(new_n331));
  INV_X1    g0131(.A(G232), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n283), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n288), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n298), .B1(G244), .B2(new_n302), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n328), .B(new_n330), .C1(new_n336), .C2(new_n312), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(new_n330), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n336), .A2(new_n305), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(G179), .C2(new_n336), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n322), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n302), .A2(G238), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n297), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(G226), .A2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n332), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n271), .C2(new_n272), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n287), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n348), .A2(KEYINPUT13), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n294), .A2(new_n296), .B1(new_n302), .B2(G238), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n288), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n346), .B(G169), .C1(new_n354), .C2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT13), .B1(new_n348), .B2(new_n353), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n358), .A3(new_n355), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(G179), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n362), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n346), .B1(new_n365), .B2(G169), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT75), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n354), .A2(new_n359), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT14), .B1(new_n368), .B2(new_n305), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT75), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n363), .A4(new_n360), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n256), .A2(G77), .ZN(new_n373));
  INV_X1    g0173(.A(G50), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n373), .B1(new_n209), .B2(G68), .C1(new_n374), .C2(new_n253), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n377), .A2(new_n378), .B1(new_n266), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT11), .B1(new_n375), .B2(new_n261), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n365), .A2(G200), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n368), .A2(G190), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(G223), .B(new_n274), .C1(new_n271), .C2(new_n272), .ZN(new_n390));
  OAI211_X1 g0190(.A(G226), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n288), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n294), .A2(new_n296), .B1(new_n302), .B2(G232), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n312), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT78), .B(new_n396), .C1(new_n397), .C2(G200), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n394), .A2(new_n395), .A3(new_n312), .ZN(new_n400));
  AOI21_X1  g0200(.A(G200), .B1(new_n394), .B2(new_n395), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n257), .A2(new_n265), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n258), .A2(new_n267), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n262), .A2(new_n264), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT77), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n266), .A2(new_n267), .A3(new_n258), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT77), .B1(new_n409), .B2(new_n404), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n201), .A2(new_n202), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G58), .A2(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n252), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n280), .A2(new_n209), .A3(new_n281), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n281), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n202), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(KEYINPUT76), .B(new_n202), .C1(new_n421), .C2(new_n422), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n423), .A2(new_n417), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n262), .B1(new_n428), .B2(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n411), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n403), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n305), .B1(new_n394), .B2(new_n395), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G179), .B2(new_n397), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT18), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT7), .B1(new_n273), .B2(new_n209), .ZN(new_n437));
  INV_X1    g0237(.A(new_n422), .ZN(new_n438));
  OAI21_X1  g0238(.A(G68), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n417), .B1(new_n439), .B2(KEYINPUT76), .ZN(new_n440));
  INV_X1    g0240(.A(new_n426), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT16), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n418), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n261), .B1(new_n443), .B2(new_n412), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n442), .A2(new_n444), .B1(new_n410), .B2(new_n408), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n397), .A2(G179), .ZN(new_n447));
  INV_X1    g0247(.A(new_n434), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n403), .A2(new_n430), .A3(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n433), .A2(new_n436), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n345), .A2(new_n385), .A3(new_n389), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT87), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n300), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n299), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(G270), .A3(new_n287), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n296), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(new_n467), .A3(G270), .A4(new_n287), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n456), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(KEYINPUT87), .A3(new_n466), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n282), .A2(G257), .A3(new_n274), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n273), .A2(G303), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n282), .A2(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(G264), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(new_n288), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n209), .C1(G33), .C2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n261), .C1(new_n209), .C2(G116), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT20), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n265), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n266), .B1(G1), .B2(new_n279), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n487), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n481), .A2(KEYINPUT21), .A3(G169), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n479), .B1(new_n470), .B2(new_n472), .ZN(new_n495));
  OAI21_X1  g0295(.A(G169), .B1(new_n486), .B2(new_n490), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(G179), .A3(new_n492), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n481), .A2(new_n312), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n491), .B1(new_n495), .B2(new_n338), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n274), .C1(new_n271), .C2(new_n272), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(KEYINPUT79), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(G1698), .B1(new_n280), .B2(new_n281), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(G244), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n506), .A2(new_n509), .A3(new_n482), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n288), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n462), .A2(G257), .A3(new_n287), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n466), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n305), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n483), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n520), .B2(new_n205), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n524));
  OAI21_X1  g0324(.A(G107), .B1(new_n437), .B2(new_n438), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n262), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n265), .A2(new_n483), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n489), .B2(new_n483), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n514), .B1(new_n511), .B2(new_n288), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(KEYINPUT82), .A3(new_n307), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT82), .B1(new_n530), .B2(new_n307), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n517), .B(new_n529), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n526), .A2(new_n528), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(G190), .ZN(new_n535));
  OAI21_X1  g0335(.A(G200), .B1(new_n530), .B2(KEYINPUT81), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n512), .A2(KEYINPUT81), .A3(new_n515), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n325), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n264), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n282), .A2(new_n209), .A3(G68), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n209), .B1(new_n352), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G87), .B2(new_n206), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n255), .B2(new_n483), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(new_n261), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT85), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  INV_X1    g0350(.A(G244), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n476), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n282), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(G238), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n283), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n287), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n460), .B(KEYINPUT83), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(G250), .A3(new_n287), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n296), .A2(new_n460), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n489), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G87), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n557), .B1(new_n552), .B2(new_n553), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(G190), .C1(new_n568), .C2(new_n287), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n549), .A2(new_n564), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n546), .A2(new_n261), .ZN(new_n571));
  INV_X1    g0371(.A(new_n540), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n548), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT85), .B(new_n540), .C1(new_n546), .C2(new_n261), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n489), .B2(new_n325), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n305), .B1(new_n559), .B2(new_n563), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n567), .B(new_n307), .C1(new_n568), .C2(new_n287), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n533), .A2(new_n538), .A3(new_n570), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n282), .A2(G257), .A3(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G294), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT90), .ZN(new_n582));
  INV_X1    g0382(.A(G250), .ZN(new_n583));
  NOR4_X1   g0383(.A1(new_n273), .A2(new_n582), .A3(new_n583), .A4(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT90), .B1(new_n507), .B2(G250), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n580), .B(new_n581), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n465), .A2(new_n288), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n288), .B1(G264), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n307), .A3(new_n466), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(G264), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n580), .A2(new_n581), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n582), .B1(new_n283), .B2(new_n583), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n507), .A2(KEYINPUT90), .A3(G250), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n466), .B(new_n590), .C1(new_n594), .C2(new_n287), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n305), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n282), .A2(new_n209), .A3(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT22), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n282), .A2(new_n599), .A3(new_n209), .A4(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n519), .A2(G20), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT23), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(KEYINPUT88), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(KEYINPUT88), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT24), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n262), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n265), .A2(new_n519), .ZN(new_n613));
  NOR2_X1   g0413(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n613), .B2(new_n614), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n565), .A2(G107), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n589), .B(new_n596), .C1(new_n612), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n588), .A2(G190), .A3(new_n466), .ZN(new_n621));
  INV_X1    g0421(.A(new_n611), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n610), .B1(new_n601), .B2(new_n607), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n261), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n595), .A2(G200), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n621), .A2(new_n624), .A3(new_n625), .A4(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n579), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n455), .A2(new_n503), .A3(new_n628), .ZN(G372));
  AND2_X1   g0429(.A1(new_n533), .A2(new_n538), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n570), .A2(new_n578), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n626), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n499), .A2(KEYINPUT91), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT91), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n493), .A2(new_n634), .A3(new_n497), .A4(new_n498), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n636), .B2(new_n620), .ZN(new_n637));
  INV_X1    g0437(.A(new_n533), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n631), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n570), .A2(new_n578), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n533), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n578), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n455), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n385), .B1(new_n388), .B2(new_n343), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n433), .A3(new_n451), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n446), .B1(new_n445), .B2(new_n449), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n435), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n450), .A2(new_n436), .A3(KEYINPUT92), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n320), .A2(new_n321), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n310), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n646), .A2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(new_n620), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT93), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n612), .B2(new_n619), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n620), .A2(new_n626), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT94), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n666), .A2(KEYINPUT94), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n664), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n491), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n503), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n636), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n499), .A2(new_n674), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n672), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT94), .B1(new_n666), .B2(new_n668), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n620), .A2(new_n664), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n686), .A3(new_n688), .ZN(G399));
  NAND2_X1  g0489(.A1(new_n212), .A2(new_n299), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n219), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n499), .A2(new_n658), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n632), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n578), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n639), .B2(new_n642), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n664), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n645), .A2(new_n674), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n567), .B1(new_n568), .B2(new_n287), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n590), .B1(new_n594), .B2(new_n287), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n706), .A3(new_n516), .ZN(new_n707));
  AOI211_X1 g0507(.A(new_n307), .B(new_n479), .C1(new_n470), .C2(new_n472), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n495), .A2(G179), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT95), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n704), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(KEYINPUT30), .A4(new_n707), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n530), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n481), .A2(new_n705), .A3(new_n595), .A4(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n664), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n628), .A2(new_n503), .A3(new_n674), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT31), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n723), .A3(new_n664), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n724), .A3(G330), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n703), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n694), .B1(new_n727), .B2(G1), .ZN(G364));
  INV_X1    g0528(.A(new_n690), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n209), .A2(G13), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n208), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n680), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n678), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n217), .B1(G20), .B2(new_n305), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n209), .A2(new_n307), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G190), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n209), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n312), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n739), .A2(new_n740), .B1(new_n743), .B2(G283), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n282), .B1(new_n747), .B2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n744), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n737), .B(KEYINPUT98), .Z(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n745), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n738), .A2(new_n312), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G326), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n312), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n307), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n757), .A2(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n755), .A2(G311), .B1(KEYINPUT100), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(KEYINPUT100), .B2(new_n764), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT101), .Z(new_n767));
  NAND2_X1  g0567(.A1(new_n753), .A2(new_n759), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n751), .B(new_n767), .C1(G322), .C2(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n282), .B1(new_n374), .B2(new_n757), .C1(new_n768), .C2(new_n201), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n746), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT99), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT32), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT32), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n762), .A2(new_n483), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G68), .B2(new_n739), .ZN(new_n778));
  INV_X1    g0578(.A(new_n750), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G87), .B1(new_n743), .B2(G107), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n771), .B(new_n781), .C1(G77), .C2(new_n755), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n736), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n678), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n736), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT97), .Z(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n212), .A2(new_n273), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n248), .A2(G45), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n300), .C2(new_n220), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n212), .A2(new_n282), .ZN(new_n796));
  INV_X1    g0596(.A(G355), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n797), .B1(G116), .B2(new_n212), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n791), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n783), .A2(new_n733), .A3(new_n788), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n735), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  OAI211_X1 g0602(.A(new_n344), .B(new_n674), .C1(new_n637), .C2(new_n644), .ZN(new_n803));
  INV_X1    g0603(.A(new_n702), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n343), .A2(new_n664), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n341), .A2(new_n664), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n337), .B2(new_n339), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n343), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n803), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n733), .B1(new_n811), .B2(new_n725), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n725), .B2(new_n811), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G137), .A2(new_n756), .B1(new_n739), .B2(G150), .ZN(new_n814));
  INV_X1    g0614(.A(G143), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n754), .B2(new_n772), .C1(new_n815), .C2(new_n768), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n282), .B1(new_n746), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G68), .B2(new_n743), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G50), .A2(new_n779), .B1(new_n761), .B2(G58), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n816), .A2(new_n817), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n273), .B1(new_n746), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n777), .B(new_n826), .C1(new_n755), .C2(G116), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n763), .B2(new_n768), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n756), .A2(G303), .B1(new_n743), .B2(G87), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n739), .A2(KEYINPUT102), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n739), .A2(KEYINPUT102), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n829), .B1(new_n519), .B2(new_n750), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n823), .A2(new_n824), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n736), .ZN(new_n836));
  INV_X1    g0636(.A(new_n733), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n736), .A2(new_n784), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n323), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n839), .C1(new_n810), .C2(new_n785), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n813), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  OR2_X1    g0642(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(G116), .A3(new_n218), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  OR3_X1    g0646(.A1(new_n219), .A2(new_n323), .A3(new_n413), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n374), .A2(G68), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n208), .B(G13), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n455), .A2(new_n722), .A3(new_n724), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT107), .Z(new_n852));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n384), .A2(new_n664), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n385), .A2(new_n389), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n384), .B(new_n664), .C1(new_n372), .C2(new_n388), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n809), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n722), .A2(new_n857), .A3(new_n724), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n428), .A2(KEYINPUT16), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n444), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n409), .A2(new_n404), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n662), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n452), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n445), .A2(new_n449), .ZN(new_n865));
  INV_X1    g0665(.A(new_n662), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n445), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n865), .A2(new_n867), .A3(new_n431), .A4(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n860), .A2(new_n861), .B1(new_n449), .B2(new_n866), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n431), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n864), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n864), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n853), .B1(new_n858), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT106), .B(new_n853), .C1(new_n858), .C2(new_n875), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(new_n867), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n430), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT17), .B1(new_n403), .B2(new_n430), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT104), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n433), .A2(new_n885), .A3(new_n451), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n652), .A2(new_n653), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT105), .B(new_n881), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n865), .A2(new_n867), .A3(new_n431), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n869), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n884), .A2(new_n886), .A3(new_n652), .A4(new_n653), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT105), .B1(new_n894), .B2(new_n881), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n880), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n873), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n858), .A2(new_n853), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n878), .A2(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(G330), .B1(new_n852), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n852), .B2(new_n901), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n385), .A2(new_n664), .ZN(new_n906));
  INV_X1    g0706(.A(new_n875), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(new_n904), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n803), .A2(new_n805), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n855), .A2(new_n856), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT103), .ZN(new_n914));
  INV_X1    g0714(.A(new_n912), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n803), .B2(new_n805), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n914), .A2(new_n918), .A3(new_n907), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n888), .A2(new_n662), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n910), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n703), .A2(new_n455), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n922), .A2(new_n656), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n903), .A2(new_n924), .B1(new_n208), .B2(new_n730), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n903), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n850), .B1(new_n925), .B2(new_n926), .ZN(G367));
  AOI21_X1  g0727(.A(new_n682), .B1(new_n671), .B2(new_n672), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n638), .A2(new_n664), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT108), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n630), .B1(new_n534), .B2(new_n674), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  INV_X1    g0734(.A(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n533), .B1(new_n935), .B2(new_n620), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n933), .A2(KEYINPUT42), .B1(new_n674), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n549), .A2(new_n566), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n664), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n631), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n697), .A2(new_n939), .A3(new_n664), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n681), .A2(new_n935), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n934), .A2(new_n937), .A3(new_n945), .A4(new_n944), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n690), .B(KEYINPUT41), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n935), .B1(new_n928), .B2(new_n687), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT44), .B(new_n935), .C1(new_n928), .C2(new_n687), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n686), .A2(new_n688), .A3(new_n932), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n688), .A4(new_n932), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n681), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n671), .A2(new_n672), .A3(new_n682), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n679), .B1(new_n969), .B2(new_n928), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n686), .A2(new_n680), .A3(new_n968), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n972), .A2(new_n726), .A3(new_n703), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n959), .A2(new_n964), .A3(new_n681), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n954), .B1(new_n975), .B2(new_n727), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n953), .B1(new_n976), .B2(new_n732), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n239), .A2(new_n792), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n789), .B1(new_n212), .B2(new_n325), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n733), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n755), .A2(G50), .B1(new_n769), .B2(G150), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n762), .A2(new_n202), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n757), .A2(new_n815), .B1(new_n201), .B2(new_n750), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G137), .C2(new_n747), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n981), .B(new_n984), .C1(new_n772), .C2(new_n832), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n742), .A2(new_n323), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n273), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT109), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n750), .A2(new_n487), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT46), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n754), .B2(new_n833), .C1(new_n749), .C2(new_n768), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n273), .B1(new_n746), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G97), .B2(new_n743), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n756), .A2(G311), .B1(new_n761), .B2(G107), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n832), .C2(new_n763), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n985), .A2(new_n988), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n980), .B1(new_n999), .B2(new_n736), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n943), .B2(new_n787), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n977), .A2(new_n1001), .ZN(G387));
  NOR2_X1   g0802(.A1(new_n973), .A2(new_n690), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n972), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n727), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n796), .A2(new_n691), .B1(G107), .B2(new_n212), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n235), .A2(new_n300), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1008));
  NOR3_X1   g0808(.A1(new_n1008), .A2(G50), .A3(new_n257), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n691), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n300), .B1(new_n202), .B2(new_n323), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1008), .B1(G50), .B2(new_n257), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n792), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1006), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n733), .B1(new_n1015), .B2(new_n790), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n673), .A2(new_n787), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n755), .A2(G303), .B1(G322), .B2(new_n756), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n825), .B2(new_n832), .C1(new_n993), .C2(new_n768), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT48), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G294), .A2(new_n779), .B1(new_n761), .B2(G283), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT49), .Z(new_n1025));
  OAI221_X1 g0825(.A(new_n273), .B1(new_n746), .B2(new_n758), .C1(new_n487), .C2(new_n742), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n768), .A2(new_n374), .B1(new_n325), .B2(new_n762), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  OAI21_X1  g0828(.A(new_n282), .B1(new_n746), .B2(new_n251), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n739), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(new_n257), .B1(new_n323), .B2(new_n750), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G97), .C2(new_n743), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n756), .A2(G159), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n755), .A2(G68), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1032), .B(new_n1035), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1025), .A2(new_n1026), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1016), .B(new_n1017), .C1(new_n736), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1004), .A2(KEYINPUT110), .A3(new_n732), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT110), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n972), .B2(new_n731), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1005), .A2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(new_n973), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n974), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n681), .B1(new_n959), .B2(new_n964), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n975), .A3(new_n729), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n789), .B1(new_n483), .B2(new_n212), .C1(new_n243), .C2(new_n792), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n282), .B1(new_n747), .B2(G322), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n519), .B2(new_n742), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n768), .A2(new_n825), .B1(new_n993), .B2(new_n757), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(G283), .C2(new_n779), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n755), .A2(G294), .B1(G116), .B2(new_n761), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n749), .B2(new_n832), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT115), .Z(new_n1057));
  NAND2_X1  g0857(.A1(new_n743), .A2(G87), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n761), .A2(G77), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n282), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n750), .A2(new_n202), .B1(new_n746), .B2(new_n815), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n832), .C2(new_n374), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1060), .B(new_n1064), .C1(new_n258), .C2(new_n755), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n768), .A2(new_n772), .B1(new_n251), .B2(new_n757), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1054), .A2(new_n1057), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n736), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n733), .B(new_n1049), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n935), .B2(new_n786), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n732), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1048), .A2(new_n1073), .ZN(G390));
  NAND3_X1  g0874(.A1(new_n726), .A2(new_n810), .A3(new_n912), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(KEYINPUT116), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n916), .A2(new_n906), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n905), .B2(new_n909), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n906), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n805), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n699), .B2(new_n808), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1084), .B2(new_n915), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n897), .B2(new_n896), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1078), .B(new_n1079), .C1(new_n1081), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT39), .B1(new_n896), .B2(new_n897), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1088), .A2(new_n908), .B1(new_n916), .B2(new_n906), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n898), .B(new_n1082), .C1(new_n915), .C2(new_n1084), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1089), .A2(new_n1077), .A3(new_n1076), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n732), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n784), .B1(new_n1088), .B2(new_n908), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n837), .B1(new_n257), .B2(new_n838), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1059), .B1(new_n768), .B2(new_n487), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT119), .Z(new_n1097));
  OAI21_X1  g0897(.A(new_n273), .B1(new_n746), .B2(new_n763), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G87), .B2(new_n779), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n756), .A2(G283), .B1(new_n743), .B2(G68), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n754), .C2(new_n483), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n832), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(G107), .B2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n819), .A2(new_n768), .B1(new_n754), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n779), .A2(G150), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n273), .B1(new_n747), .B2(G125), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n374), .B2(new_n742), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n756), .A2(G128), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n772), .B2(new_n762), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n1102), .C2(G137), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1097), .A2(new_n1103), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1094), .B(new_n1095), .C1(new_n1069), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n455), .A2(new_n726), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n922), .A2(new_n656), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n915), .B1(new_n725), .B2(new_n809), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1075), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n911), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1075), .A2(new_n1084), .A3(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n690), .B1(new_n1128), .B2(new_n1092), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1087), .A3(new_n1127), .A4(new_n1091), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1118), .A2(new_n1131), .ZN(G378));
  INV_X1    g0932(.A(new_n1120), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1092), .B2(new_n1125), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n910), .A2(new_n919), .A3(new_n920), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT122), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n270), .A2(new_n662), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n322), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n322), .A2(new_n1138), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n322), .A2(new_n1138), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n1139), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1136), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1143), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT122), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n878), .A2(new_n879), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n898), .A2(new_n899), .ZN(new_n1153));
  AND4_X1   g0953(.A1(G330), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n900), .B2(G330), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1135), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(G330), .A3(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1155), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n900), .A2(G330), .A3(new_n1151), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n921), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1134), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT57), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1125), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1158), .B(new_n1162), .C1(new_n1167), .C2(new_n1133), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n729), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1158), .A2(new_n732), .A3(new_n1162), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n838), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n733), .B1(G50), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT121), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n982), .B1(G283), .B2(new_n747), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n325), .B2(new_n754), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n742), .A2(new_n201), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1030), .A2(new_n483), .B1(new_n757), .B2(new_n487), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n273), .A2(new_n299), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n779), .B2(G77), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1179), .C1(KEYINPUT120), .C2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1181), .A2(KEYINPUT120), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1177), .B(new_n1184), .C1(G107), .C2(new_n769), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  INV_X1    g0987(.A(G137), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1187), .A2(new_n768), .B1(new_n754), .B2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n756), .A2(G125), .B1(new_n761), .B2(G150), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n819), .B2(new_n1030), .C1(new_n750), .C2(new_n1104), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n743), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1180), .B(new_n374), .C1(G33), .C2(G41), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n1186), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1175), .B1(new_n1069), .B2(new_n1201), .C1(new_n1151), .C2(new_n785), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1172), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1171), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n1133), .A2(new_n1166), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n954), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1126), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n733), .B1(G68), .B2(new_n1173), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n755), .A2(G107), .B1(new_n769), .B2(G283), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n761), .A2(new_n539), .B1(new_n747), .B2(G303), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n756), .A2(G294), .B1(new_n779), .B2(G97), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT123), .B1(new_n986), .B2(new_n282), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n986), .A2(KEYINPUT123), .A3(new_n282), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n832), .C2(new_n487), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n273), .B(new_n1178), .C1(G128), .C2(new_n747), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n754), .B2(new_n251), .C1(new_n1188), .C2(new_n768), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G159), .A2(new_n779), .B1(new_n761), .B2(G50), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n819), .B2(new_n757), .C1(new_n832), .C2(new_n1104), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1213), .A2(new_n1216), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1209), .B1(new_n1221), .B2(new_n736), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n912), .B2(new_n785), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1166), .B2(new_n731), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1208), .A2(new_n1225), .ZN(G381));
  XNOR2_X1  g1026(.A(G375), .B(KEYINPUT124), .ZN(new_n1227));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n841), .A3(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1230), .A2(G387), .A3(G381), .ZN(new_n1231));
  OR3_X1    g1031(.A1(new_n1227), .A2(G378), .A3(new_n1231), .ZN(G407));
  NAND2_X1  g1032(.A1(new_n663), .A2(G213), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n1227), .A2(G378), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(new_n1234), .A3(G213), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1203), .B1(new_n1164), .B2(new_n1207), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(G378), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n729), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1092), .A2(new_n1125), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1120), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G378), .B(new_n1204), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1117), .B1(new_n1130), .B2(new_n1129), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1168), .A2(new_n954), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(KEYINPUT125), .C1(new_n1246), .C2(new_n1203), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1238), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1133), .A2(new_n1166), .A3(KEYINPUT60), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1249), .A2(new_n729), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1206), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n841), .B1(new_n1253), .B2(new_n1224), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1225), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1248), .A2(new_n1233), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT126), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1248), .A2(new_n1233), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1254), .A2(new_n1256), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1248), .A2(new_n1233), .A3(new_n1258), .A4(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1262), .A2(new_n1268), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n977), .A2(new_n1001), .A3(G390), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G390), .B1(new_n977), .B2(new_n1001), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n801), .B1(new_n1005), .B2(new_n1042), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1273), .A2(new_n1274), .B1(new_n1229), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1228), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1229), .A2(new_n1275), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n977), .A2(G390), .A3(new_n1001), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n1259), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1284), .B(new_n1285), .C1(new_n1283), .C2(new_n1259), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1245), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1257), .A3(new_n1244), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G378), .B1(new_n1171), .B2(new_n1204), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1244), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1258), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1281), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1281), .B1(new_n1292), .B2(new_n1289), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI211_X1 g1096(.A(KEYINPUT127), .B(new_n1281), .C1(new_n1292), .C2(new_n1289), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


