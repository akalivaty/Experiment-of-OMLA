//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  AND2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(KEYINPUT14), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT15), .A4(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT15), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT14), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n217), .A2(new_n212), .A3(KEYINPUT15), .A4(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n213), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT93), .ZN(new_n223));
  INV_X1    g022(.A(G8gat), .ZN(new_n224));
  INV_X1    g023(.A(G22gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G15gat), .ZN(new_n226));
  INV_X1    g025(.A(G15gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G22gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT94), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT94), .B1(new_n226), .B2(new_n228), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G1gat), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n228), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(G1gat), .B1(new_n237), .B2(new_n229), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT95), .B(new_n224), .C1(new_n234), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT93), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(new_n213), .C1(new_n214), .C2(new_n221), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n237), .B(new_n229), .C1(new_n232), .C2(G1gat), .ZN(new_n242));
  INV_X1    g041(.A(G1gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n230), .B2(new_n231), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(KEYINPUT95), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n224), .A2(KEYINPUT95), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n223), .A2(new_n239), .A3(new_n241), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  INV_X1    g049(.A(new_n241), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n217), .A2(new_n212), .A3(new_n218), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n219), .A3(new_n220), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n240), .B1(new_n255), .B2(new_n213), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n247), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n249), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G229gat), .A2(G233gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT18), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(G229gat), .B2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n223), .A2(new_n241), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(new_n250), .ZN(new_n268));
  INV_X1    g067(.A(new_n260), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n248), .B(new_n265), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n262), .B(KEYINPUT13), .Z(new_n271));
  AOI22_X1  g070(.A1(new_n223), .A2(new_n241), .B1(new_n239), .B2(new_n247), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n249), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n206), .B1(new_n263), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n260), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(new_n248), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n261), .B2(new_n265), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n262), .B(new_n248), .C1(new_n268), .C2(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n264), .ZN(new_n281));
  INV_X1    g080(.A(new_n206), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G127gat), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G134gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n293), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT1), .B1(new_n287), .B2(new_n291), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n294), .A3(G127gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT68), .B1(new_n294), .B2(G127gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n296), .A2(G134gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT69), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n300), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI211_X1 g110(.A(KEYINPUT70), .B(new_n300), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n299), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G141gat), .B(G148gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G141gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n320), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n320), .A2(new_n328), .A3(KEYINPUT83), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT83), .B1(new_n320), .B2(new_n328), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n334), .B2(KEYINPUT3), .ZN(new_n335));
  NOR4_X1   g134(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT84), .A4(new_n329), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n313), .B(new_n330), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n320), .A2(new_n328), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(new_n299), .C1(new_n311), .C2(new_n312), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n299), .ZN(new_n342));
  INV_X1    g141(.A(new_n308), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n295), .A2(new_n297), .A3(KEYINPUT68), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT69), .B1(new_n344), .B2(new_n302), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT70), .B1(new_n346), .B2(new_n300), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n309), .A2(new_n310), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n337), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n313), .A2(new_n334), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n354), .B2(new_n339), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  OAI22_X1  g155(.A1(new_n351), .A2(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n350), .A2(new_n341), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n358), .A2(KEYINPUT5), .A3(new_n352), .A4(new_n337), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT85), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(new_n359), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n363), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n357), .A2(new_n359), .A3(new_n370), .A4(new_n364), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(new_n368), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n365), .A2(new_n369), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  XOR2_X1   g173(.A(G211gat), .B(G218gat), .Z(new_n375));
  INV_X1    g174(.A(G197gat), .ZN(new_n376));
  INV_X1    g175(.A(G204gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  NAND2_X1  g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n378), .A2(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n380), .ZN(new_n385));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386));
  AND2_X1   g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n374), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n388), .B2(new_n375), .ZN(new_n392));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(KEYINPUT81), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n388), .B2(KEYINPUT79), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n382), .A2(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT80), .A3(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n390), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  INV_X1    g199(.A(G169gat), .ZN(new_n401));
  INV_X1    g200(.A(G176gat), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n400), .A2(KEYINPUT24), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G183gat), .ZN(new_n405));
  INV_X1    g204(.A(G190gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT24), .A3(new_n400), .ZN(new_n408));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n404), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n404), .A2(new_n413), .A3(KEYINPUT25), .A4(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n420));
  OR3_X1    g219(.A1(new_n419), .A2(new_n409), .A3(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(KEYINPUT66), .A2(KEYINPUT26), .ZN(new_n422));
  NAND2_X1  g221(.A1(KEYINPUT66), .A2(KEYINPUT26), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n419), .B2(new_n409), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n405), .A2(KEYINPUT27), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G183gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n429), .A3(new_n406), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n426), .B(new_n400), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n418), .B1(new_n436), .B2(KEYINPUT67), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(KEYINPUT67), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n418), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n439), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n399), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT28), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n433), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n426), .A4(new_n400), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(new_n418), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n440), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n443), .A2(new_n440), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT82), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n400), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n448), .B2(new_n433), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n458), .B2(new_n426), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n444), .B1(new_n437), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n439), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n446), .B1(new_n464), .B2(new_n399), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n390), .A2(new_n395), .A3(new_n398), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n456), .B2(new_n463), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n446), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(new_n475), .A3(new_n468), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n372), .A2(new_n373), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n438), .A2(new_n349), .A3(KEYINPUT73), .A4(new_n441), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n452), .B2(new_n313), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n452), .A2(new_n313), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n485), .ZN(new_n488));
  XOR2_X1   g287(.A(KEYINPUT74), .B(KEYINPUT33), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT75), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G71gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(G99gat), .Z(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n481), .A3(new_n484), .A4(new_n482), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT77), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT34), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT34), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n489), .B1(new_n483), .B2(new_n485), .ZN(new_n502));
  INV_X1    g301(.A(new_n495), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n486), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT78), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n496), .A2(new_n501), .A3(new_n507), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G50gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  INV_X1    g312(.A(new_n334), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n471), .A2(new_n444), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(new_n329), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n330), .A2(new_n444), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n390), .A3(new_n395), .A4(new_n398), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(G228gat), .A3(G233gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n513), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n399), .B2(new_n517), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT3), .B1(new_n471), .B2(new_n444), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(KEYINPUT88), .C1(new_n514), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n521), .B(KEYINPUT86), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n395), .A2(KEYINPUT87), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n392), .A2(new_n529), .A3(new_n394), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n382), .B2(new_n393), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n444), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n338), .B1(new_n532), .B2(new_n329), .ZN(new_n533));
  INV_X1    g332(.A(new_n518), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n512), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(G22gat), .B1(new_n536), .B2(KEYINPUT89), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n527), .B(new_n530), .C1(new_n382), .C2(new_n393), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT3), .B1(new_n538), .B2(new_n444), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n518), .B1(new_n539), .B2(new_n338), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n520), .A2(new_n524), .B1(new_n540), .B2(new_n526), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(new_n512), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n543), .B(new_n225), .C1(new_n541), .C2(new_n512), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n537), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n537), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n486), .A2(new_n502), .A3(new_n503), .ZN(new_n548));
  AOI221_X4 g347(.A(new_n478), .B1(new_n495), .B2(new_n489), .C1(new_n483), .C2(new_n485), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT76), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n501), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n496), .A2(new_n552), .A3(new_n504), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n477), .A2(new_n509), .A3(new_n547), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n501), .B1(new_n496), .B2(new_n504), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n506), .B2(new_n508), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT35), .B1(new_n474), .B2(new_n476), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n365), .A2(KEYINPUT92), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n357), .A2(new_n359), .A3(new_n561), .A4(new_n364), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n560), .A2(new_n368), .A3(new_n369), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n373), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n558), .A2(new_n559), .A3(new_n547), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n509), .A2(new_n554), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n568));
  INV_X1    g367(.A(new_n446), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT82), .B1(new_n460), .B2(new_n439), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n461), .A2(new_n454), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(KEYINPUT82), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(new_n471), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n470), .B1(new_n573), .B2(KEYINPUT37), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n465), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT38), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n468), .B1(new_n465), .B2(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n464), .A2(new_n471), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n442), .A2(new_n445), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n580), .B2(new_n399), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT38), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n578), .A2(new_n582), .B1(new_n465), .B2(new_n468), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n577), .A2(new_n583), .A3(new_n373), .A4(new_n563), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n351), .A2(new_n353), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n363), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n354), .A2(new_n352), .A3(new_n339), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT39), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n353), .B2(new_n351), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(KEYINPUT91), .B(new_n585), .C1(new_n588), .C2(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n351), .A2(new_n353), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT39), .A3(new_n589), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(KEYINPUT40), .A3(new_n363), .A4(new_n587), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n560), .A2(new_n599), .A3(new_n562), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n596), .A2(new_n600), .A3(new_n476), .A4(new_n474), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n601), .A3(new_n547), .ZN(new_n602));
  INV_X1    g401(.A(new_n547), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n372), .A2(new_n373), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n474), .A2(new_n476), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n558), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n568), .A2(new_n602), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n285), .B1(new_n566), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT97), .A3(new_n615), .ZN(new_n619));
  INV_X1    g418(.A(G57gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G64gat), .ZN(new_n621));
  INV_X1    g420(.A(G64gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G57gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n614), .ZN(new_n627));
  NOR3_X1   g426(.A1(KEYINPUT96), .A2(G71gat), .A3(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT98), .B1(new_n622), .B2(G57gat), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n620), .A3(G64gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n633), .A3(new_n623), .ZN(new_n634));
  XNOR2_X1  g433(.A(G71gat), .B(G78gat), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n619), .A4(new_n618), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT20), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(new_n640), .ZN(new_n646));
  INV_X1    g445(.A(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n613), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n260), .B1(new_n638), .B2(new_n637), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(new_n648), .A3(new_n613), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n653), .B1(new_n657), .B2(new_n649), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G99gat), .B(G106gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G85gat), .A2(G92gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT100), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(G85gat), .A3(G92gat), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT7), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT7), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(KEYINPUT100), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  INV_X1    g468(.A(G92gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G99gat), .A2(G106gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT8), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n661), .B1(new_n666), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT7), .ZN(new_n676));
  AOI22_X1  g475(.A1(KEYINPUT8), .A2(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n660), .A3(new_n668), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n259), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n223), .A2(new_n241), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT101), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(G190gat), .B(G218gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n680), .B(new_n689), .C1(new_n684), .C2(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G134gat), .B(G162gat), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n688), .B(new_n690), .C1(new_n698), .C2(new_n695), .ZN(new_n699));
  INV_X1    g498(.A(G230gat), .ZN(new_n700));
  INV_X1    g499(.A(G233gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n678), .B(new_n675), .C1(new_n637), .C2(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n618), .A2(new_n635), .A3(new_n619), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n706), .A2(new_n634), .B1(new_n625), .B2(new_n629), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n678), .A2(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n679), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT10), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT10), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n679), .A2(new_n637), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n703), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n705), .A2(new_n702), .A3(new_n709), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(G120gat), .B(G148gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(G176gat), .B(G204gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n716), .B(new_n717), .Z(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n714), .A2(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n714), .A2(KEYINPUT104), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n721), .A2(new_n713), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n659), .A2(new_n697), .A3(new_n699), .A4(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n611), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n604), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n243), .ZN(G1324gat));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n605), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT16), .B(G8gat), .Z(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G8gat), .B1(new_n728), .B2(new_n605), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n736));
  MUX2_X1   g535(.A(KEYINPUT105), .B(new_n736), .S(new_n733), .Z(new_n737));
  AOI22_X1  g536(.A1(new_n734), .A2(new_n735), .B1(new_n732), .B2(new_n737), .ZN(G1325gat));
  AOI21_X1  g537(.A(new_n608), .B1(new_n509), .B2(new_n554), .ZN(new_n739));
  AOI211_X1 g538(.A(KEYINPUT36), .B(new_n557), .C1(new_n506), .C2(new_n508), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G15gat), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n558), .A2(new_n227), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n728), .B2(new_n743), .ZN(G1326gat));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n547), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT43), .B(G22gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1327gat));
  INV_X1    g546(.A(new_n659), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n725), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n697), .A2(new_n699), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n611), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(G29gat), .A3(new_n604), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT45), .Z(new_n755));
  INV_X1    g554(.A(new_n604), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n275), .A2(KEYINPUT106), .A3(new_n283), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT106), .B1(new_n275), .B2(new_n283), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n749), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n566), .A2(new_n610), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n750), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n750), .A2(new_n761), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT107), .B1(new_n477), .B2(new_n547), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n603), .A2(new_n606), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n741), .A2(new_n602), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(new_n768), .B2(new_n566), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n756), .B(new_n760), .C1(new_n763), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n215), .B1(new_n770), .B2(KEYINPUT108), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT108), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n772), .ZN(G1328gat));
  NOR3_X1   g572(.A1(new_n753), .A2(G36gat), .A3(new_n605), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT46), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n763), .A2(new_n769), .ZN(new_n776));
  INV_X1    g575(.A(new_n605), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n760), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n216), .B2(new_n779), .ZN(G1329gat));
  NAND2_X1  g579(.A1(new_n568), .A2(new_n609), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(new_n760), .C1(new_n763), .C2(new_n769), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G43gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n558), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n753), .A2(G43gat), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n783), .B2(new_n785), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1330gat));
  INV_X1    g588(.A(G50gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n547), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n760), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n753), .B2(new_n547), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT48), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1331gat));
  NAND3_X1  g597(.A1(new_n568), .A2(new_n602), .A3(new_n609), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n767), .A2(new_n765), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n566), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n263), .A2(new_n274), .A3(new_n206), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n282), .B1(new_n279), .B2(new_n281), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n275), .A2(KEYINPUT106), .A3(new_n283), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR4_X1   g606(.A1(new_n807), .A2(new_n748), .A3(new_n750), .A4(new_n725), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n604), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(new_n620), .ZN(G1332gat));
  AND3_X1   g610(.A1(new_n801), .A2(KEYINPUT109), .A3(new_n808), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT109), .B1(new_n801), .B2(new_n808), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n605), .ZN(new_n814));
  NOR2_X1   g613(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n815));
  AND2_X1   g614(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n814), .B2(new_n815), .ZN(G1333gat));
  NOR3_X1   g617(.A1(new_n812), .A2(new_n813), .A3(new_n741), .ZN(new_n819));
  INV_X1    g618(.A(G71gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n558), .A2(new_n820), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n819), .A2(new_n820), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI221_X1 g623(.A(KEYINPUT50), .B1(new_n809), .B2(new_n821), .C1(new_n819), .C2(new_n820), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1334gat));
  NOR3_X1   g625(.A1(new_n812), .A2(new_n813), .A3(new_n547), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g627(.A1(new_n807), .A2(new_n659), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT110), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n725), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n776), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G85gat), .B1(new_n832), .B2(new_n604), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n830), .A2(new_n751), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n801), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n801), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n724), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n756), .A2(new_n669), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  OAI211_X1 g638(.A(new_n777), .B(new_n831), .C1(new_n763), .C2(new_n769), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G92gat), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n605), .A2(G92gat), .A3(new_n725), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT112), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n835), .B2(new_n836), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n841), .B(new_n844), .C1(new_n847), .C2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1337gat));
  OAI21_X1  g650(.A(G99gat), .B1(new_n832), .B2(new_n741), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n784), .A2(G99gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n837), .B2(new_n853), .ZN(G1338gat));
  OAI211_X1 g653(.A(new_n603), .B(new_n831), .C1(new_n763), .C2(new_n769), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G106gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n547), .A2(G106gat), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n724), .B(new_n857), .C1(new_n835), .C2(new_n836), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1339gat));
  NAND3_X1  g662(.A1(new_n727), .A2(new_n759), .A3(KEYINPUT114), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n807), .B2(new_n726), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n723), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n869), .B(new_n703), .C1(new_n710), .C2(new_n712), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n719), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(KEYINPUT115), .A3(new_n719), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n707), .A2(new_n679), .A3(new_n708), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n679), .B1(new_n707), .B2(new_n708), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n711), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n712), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n702), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n880), .A2(new_n713), .A3(KEYINPUT54), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n868), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n713), .A3(KEYINPUT54), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n870), .A2(KEYINPUT115), .A3(new_n719), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT115), .B1(new_n870), .B2(new_n719), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n882), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n261), .A2(new_n262), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n249), .A2(new_n272), .A3(new_n271), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n205), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n283), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n890), .A2(new_n750), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n283), .A2(new_n893), .A3(new_n724), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n890), .B2(new_n807), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n750), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n867), .B1(new_n898), .B2(new_n748), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n604), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n567), .A2(new_n603), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n605), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT116), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n290), .A3(new_n807), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n899), .A2(new_n603), .A3(new_n784), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n777), .A2(new_n604), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G113gat), .B1(new_n907), .B2(new_n285), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n904), .A2(new_n908), .ZN(G1340gat));
  NAND3_X1  g708(.A1(new_n903), .A2(new_n286), .A3(new_n724), .ZN(new_n910));
  OAI21_X1  g709(.A(G120gat), .B1(new_n907), .B2(new_n725), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1341gat));
  OAI21_X1  g711(.A(G127gat), .B1(new_n907), .B2(new_n748), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n659), .A2(new_n296), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n902), .B2(new_n914), .ZN(G1342gat));
  OR3_X1    g714(.A1(new_n902), .A2(G134gat), .A3(new_n751), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n917));
  OAI21_X1  g716(.A(G134gat), .B1(new_n907), .B2(new_n751), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G1343gat));
  NOR2_X1   g719(.A1(new_n781), .A2(new_n547), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT120), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n900), .A2(new_n605), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n285), .A2(G141gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n603), .A2(KEYINPUT57), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n881), .B1(new_n873), .B2(new_n874), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT118), .B1(new_n928), .B2(KEYINPUT55), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n888), .A2(new_n930), .A3(new_n882), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n929), .A2(new_n284), .A3(new_n884), .A4(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n896), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n751), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n659), .B1(new_n935), .B2(new_n895), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n927), .B1(new_n936), .B2(new_n867), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n884), .B(new_n889), .C1(new_n757), .C2(new_n758), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n750), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n890), .A2(new_n750), .A3(new_n894), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n748), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n867), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n547), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n937), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n741), .A2(new_n906), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n284), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G141gat), .ZN(new_n950));
  XOR2_X1   g749(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n951));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n946), .B2(new_n948), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n946), .A2(new_n953), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n807), .A3(new_n956), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n957), .A2(G141gat), .B1(new_n924), .B2(new_n925), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT58), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(G1344gat));
  INV_X1    g759(.A(KEYINPUT59), .ZN(new_n961));
  AOI211_X1 g760(.A(new_n961), .B(G148gat), .C1(new_n924), .C2(new_n724), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n945), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n726), .A2(new_n284), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n936), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n547), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n966), .B2(KEYINPUT57), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n725), .A2(new_n961), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n967), .A2(new_n741), .A3(new_n906), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n944), .B1(new_n899), .B2(new_n547), .ZN(new_n970));
  AOI211_X1 g769(.A(KEYINPUT119), .B(new_n947), .C1(new_n970), .C2(new_n937), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n971), .A2(new_n954), .A3(new_n725), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(KEYINPUT59), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n962), .B1(new_n973), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g773(.A(G155gat), .B1(new_n924), .B2(new_n659), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n971), .A2(new_n954), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n659), .A2(G155gat), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT122), .Z(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n976), .B2(new_n978), .ZN(G1346gat));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n980));
  INV_X1    g779(.A(G162gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n981), .B1(new_n976), .B2(new_n750), .ZN(new_n982));
  NOR4_X1   g781(.A1(new_n922), .A2(G162gat), .A3(new_n923), .A4(new_n751), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n924), .A2(new_n981), .A3(new_n750), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n971), .A2(new_n954), .A3(new_n751), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n985), .B(KEYINPUT123), .C1(new_n981), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n987), .ZN(G1347gat));
  NOR2_X1   g787(.A1(new_n756), .A2(new_n605), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n905), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n990), .A2(new_n401), .A3(new_n285), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n899), .A2(new_n756), .A3(new_n605), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(new_n901), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n807), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n991), .B1(new_n401), .B2(new_n995), .ZN(G1348gat));
  OAI21_X1  g795(.A(G176gat), .B1(new_n990), .B2(new_n725), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n724), .A2(new_n402), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n993), .B2(new_n998), .ZN(G1349gat));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n1000), .B1(new_n990), .B2(new_n748), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n905), .A2(KEYINPUT124), .A3(new_n659), .A4(new_n989), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1001), .A2(G183gat), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n994), .A2(new_n427), .A3(new_n429), .A4(new_n659), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g805(.A1(new_n994), .A2(new_n406), .A3(new_n750), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n905), .A2(new_n750), .A3(new_n989), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n1010));
  AND4_X1   g809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(G190gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n406), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n1012));
  AOI22_X1  g811(.A1(new_n1009), .A2(new_n1012), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1007), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1016));
  OAI211_X1 g815(.A(new_n1016), .B(new_n1007), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1015), .A2(new_n1017), .ZN(G1351gat));
  NAND3_X1  g817(.A1(new_n967), .A2(new_n741), .A3(new_n989), .ZN(new_n1019));
  NOR3_X1   g818(.A1(new_n1019), .A2(new_n376), .A3(new_n285), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n992), .A2(new_n921), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g821(.A(G197gat), .B1(new_n1022), .B2(new_n807), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n1020), .A2(new_n1023), .ZN(G1352gat));
  XNOR2_X1  g823(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1025));
  NOR3_X1   g824(.A1(new_n1021), .A2(new_n725), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1025), .B1(new_n1019), .B2(new_n725), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(new_n1028), .ZN(G1353gat));
  OR3_X1    g828(.A1(new_n1021), .A2(G211gat), .A3(new_n748), .ZN(new_n1030));
  NAND4_X1  g829(.A1(new_n967), .A2(new_n741), .A3(new_n659), .A4(new_n989), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1031), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(KEYINPUT63), .B1(new_n1031), .B2(G211gat), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(G1354gat));
  OAI21_X1  g833(.A(G218gat), .B1(new_n1019), .B2(new_n751), .ZN(new_n1035));
  OR2_X1    g834(.A1(new_n751), .A2(G218gat), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1035), .B1(new_n1021), .B2(new_n1036), .ZN(G1355gat));
endmodule


