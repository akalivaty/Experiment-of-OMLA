

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592;

  INV_X1 U327 ( .A(n574), .ZN(n383) );
  AND2_X1 U328 ( .A1(n384), .A2(n383), .ZN(n295) );
  XOR2_X1 U329 ( .A(KEYINPUT89), .B(G218GAT), .Z(n296) );
  XOR2_X1 U330 ( .A(KEYINPUT58), .B(n571), .Z(n297) );
  AND2_X1 U331 ( .A1(n507), .A2(n506), .ZN(n508) );
  INV_X1 U332 ( .A(KEYINPUT23), .ZN(n357) );
  XNOR2_X1 U333 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U334 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U335 ( .A(KEYINPUT48), .B(n516), .ZN(n549) );
  INV_X1 U336 ( .A(n589), .ZN(n470) );
  OR2_X1 U337 ( .A1(n575), .A2(n554), .ZN(n555) );
  NAND2_X1 U338 ( .A1(n470), .A2(n566), .ZN(n471) );
  OR2_X1 U339 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U340 ( .A(n372), .B(n371), .Z(n552) );
  XNOR2_X1 U341 ( .A(n461), .B(n460), .ZN(n581) );
  XOR2_X1 U342 ( .A(KEYINPUT38), .B(n475), .Z(n483) );
  XNOR2_X1 U343 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n463) );
  XOR2_X1 U344 ( .A(G57GAT), .B(G120GAT), .Z(n299) );
  XNOR2_X1 U345 ( .A(G141GAT), .B(G1GAT), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U347 ( .A(G85GAT), .B(G148GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n320) );
  XOR2_X1 U351 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT4), .B(KEYINPUT98), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U357 ( .A(n309), .B(n308), .Z(n318) );
  XOR2_X1 U358 ( .A(KEYINPUT90), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(n312), .Z(n368) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n313), .B(G127GAT), .ZN(n328) );
  XOR2_X1 U364 ( .A(n328), .B(KEYINPUT94), .Z(n315) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n368), .B(n316), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n574) );
  XOR2_X1 U370 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n322) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G15GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n338) );
  XOR2_X1 U373 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n324) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n325), .B(KEYINPUT20), .Z(n330) );
  XOR2_X1 U377 ( .A(G183GAT), .B(KEYINPUT17), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n345) );
  XNOR2_X1 U380 ( .A(n328), .B(n345), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U382 ( .A(G176GAT), .B(KEYINPUT80), .Z(n332) );
  XOR2_X1 U383 ( .A(G190GAT), .B(G134GAT), .Z(n420) );
  XOR2_X1 U384 ( .A(G120GAT), .B(G71GAT), .Z(n459) );
  XNOR2_X1 U385 ( .A(n420), .B(n459), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U387 ( .A(n334), .B(n333), .Z(n336) );
  XNOR2_X1 U388 ( .A(G43GAT), .B(G99GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X2 U390 ( .A(n338), .B(n337), .Z(n556) );
  XOR2_X1 U391 ( .A(KEYINPUT74), .B(G204GAT), .Z(n340) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G190GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n349) );
  XOR2_X1 U394 ( .A(G169GAT), .B(G8GAT), .Z(n438) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n341), .B(G64GAT), .ZN(n443) );
  XOR2_X1 U397 ( .A(n438), .B(n443), .Z(n343) );
  NAND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U400 ( .A(n344), .B(KEYINPUT100), .Z(n347) );
  XNOR2_X1 U401 ( .A(n345), .B(KEYINPUT99), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n352) );
  XNOR2_X1 U404 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n296), .B(n350), .ZN(n351) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(n351), .ZN(n360) );
  XNOR2_X1 U407 ( .A(n352), .B(n360), .ZN(n548) );
  XNOR2_X1 U408 ( .A(KEYINPUT27), .B(n548), .ZN(n379) );
  NAND2_X1 U409 ( .A1(n574), .A2(n379), .ZN(n517) );
  NOR2_X1 U410 ( .A1(n556), .A2(n517), .ZN(n373) );
  XOR2_X1 U411 ( .A(G78GAT), .B(G148GAT), .Z(n354) );
  XNOR2_X1 U412 ( .A(G106GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n451) );
  XOR2_X1 U414 ( .A(n451), .B(KEYINPUT93), .Z(n356) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n372) );
  XOR2_X1 U417 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n358) );
  XOR2_X1 U418 ( .A(n361), .B(KEYINPUT85), .Z(n370) );
  XOR2_X1 U419 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n363) );
  XNOR2_X1 U420 ( .A(KEYINPUT91), .B(KEYINPUT88), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U422 ( .A(n364), .B(KEYINPUT92), .Z(n366) );
  XOR2_X1 U423 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(n439), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n552), .B(KEYINPUT28), .ZN(n520) );
  NAND2_X1 U429 ( .A1(n373), .A2(n520), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(KEYINPUT101), .ZN(n385) );
  NAND2_X1 U431 ( .A1(n556), .A2(n548), .ZN(n375) );
  XNOR2_X1 U432 ( .A(KEYINPUT102), .B(n375), .ZN(n376) );
  NAND2_X1 U433 ( .A1(n376), .A2(n552), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n377), .B(KEYINPUT25), .ZN(n381) );
  NOR2_X1 U435 ( .A1(n556), .A2(n552), .ZN(n378) );
  XNOR2_X1 U436 ( .A(KEYINPUT26), .B(n378), .ZN(n577) );
  AND2_X1 U437 ( .A1(n379), .A2(n577), .ZN(n380) );
  NOR2_X1 U438 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT103), .ZN(n384) );
  NOR2_X1 U440 ( .A1(n385), .A2(n295), .ZN(n472) );
  XOR2_X1 U441 ( .A(KEYINPUT13), .B(G57GAT), .Z(n458) );
  XOR2_X1 U442 ( .A(G211GAT), .B(G78GAT), .Z(n387) );
  XNOR2_X1 U443 ( .A(G22GAT), .B(G155GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U445 ( .A(n458), .B(n388), .Z(n390) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n391), .B(KEYINPUT12), .Z(n394) );
  XNOR2_X1 U449 ( .A(G15GAT), .B(G1GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT67), .ZN(n436) );
  XNOR2_X1 U451 ( .A(n436), .B(KEYINPUT79), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT74), .B(G71GAT), .Z(n396) );
  XNOR2_X1 U454 ( .A(G127GAT), .B(G183GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U456 ( .A(n398), .B(n397), .Z(n406) );
  XOR2_X1 U457 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n402) );
  XNOR2_X1 U461 ( .A(G8GAT), .B(G64GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n566) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n407), .B(G29GAT), .ZN(n408) );
  XOR2_X1 U467 ( .A(n408), .B(KEYINPUT8), .Z(n410) );
  XNOR2_X1 U468 ( .A(G43GAT), .B(G50GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n433) );
  XOR2_X1 U470 ( .A(G99GAT), .B(G85GAT), .Z(n442) );
  XOR2_X1 U471 ( .A(KEYINPUT73), .B(n442), .Z(n412) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U474 ( .A(KEYINPUT10), .B(G92GAT), .Z(n414) );
  XNOR2_X1 U475 ( .A(G162GAT), .B(G106GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U477 ( .A(n416), .B(n415), .Z(n422) );
  XOR2_X1 U478 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n418) );
  XNOR2_X1 U479 ( .A(G218GAT), .B(KEYINPUT72), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n433), .B(n423), .ZN(n546) );
  NOR2_X1 U484 ( .A1(n566), .A2(n546), .ZN(n424) );
  XOR2_X1 U485 ( .A(KEYINPUT16), .B(n424), .Z(n425) );
  NOR2_X1 U486 ( .A1(n472), .A2(n425), .ZN(n426) );
  XOR2_X1 U487 ( .A(KEYINPUT104), .B(n426), .Z(n485) );
  XOR2_X1 U488 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n428) );
  NAND2_X1 U489 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U491 ( .A(n429), .B(KEYINPUT66), .Z(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n431) );
  XNOR2_X1 U493 ( .A(G197GAT), .B(G113GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U497 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n578) );
  XOR2_X1 U500 ( .A(n578), .B(KEYINPUT68), .Z(n558) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n445) );
  AND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n448) );
  INV_X1 U504 ( .A(n448), .ZN(n446) );
  NAND2_X1 U505 ( .A1(n446), .A2(KEYINPUT33), .ZN(n450) );
  INV_X1 U506 ( .A(KEYINPUT33), .ZN(n447) );
  NAND2_X1 U507 ( .A1(n448), .A2(n447), .ZN(n449) );
  NAND2_X1 U508 ( .A1(n450), .A2(n449), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n451), .B(KEYINPUT32), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n454) );
  XOR2_X1 U513 ( .A(n455), .B(n454), .Z(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(n460) );
  OR2_X1 U516 ( .A1(n558), .A2(n581), .ZN(n474) );
  NOR2_X1 U517 ( .A1(n485), .A2(n474), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n574), .A2(n468), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(G1324GAT) );
  NAND2_X1 U520 ( .A1(n548), .A2(n468), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U522 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n466) );
  NAND2_X1 U523 ( .A1(n468), .A2(n556), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U525 ( .A(G15GAT), .B(n467), .Z(G1326GAT) );
  INV_X1 U526 ( .A(n520), .ZN(n501) );
  NAND2_X1 U527 ( .A1(n468), .A2(n501), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U529 ( .A(G29GAT), .B(KEYINPUT39), .Z(n477) );
  INV_X1 U530 ( .A(n546), .ZN(n570) );
  XNOR2_X1 U531 ( .A(n570), .B(KEYINPUT36), .ZN(n589) );
  XOR2_X1 U532 ( .A(KEYINPUT37), .B(n473), .Z(n495) );
  OR2_X1 U533 ( .A1(n495), .A2(n474), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n574), .A2(n483), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(G1328GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n479) );
  NAND2_X1 U537 ( .A1(n483), .A2(n548), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G36GAT), .B(n480), .ZN(G1329GAT) );
  NAND2_X1 U540 ( .A1(n483), .A2(n556), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT40), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G43GAT), .B(n482), .ZN(G1330GAT) );
  NAND2_X1 U543 ( .A1(n501), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(G50GAT), .B(n484), .ZN(G1331GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT41), .B(n581), .Z(n540) );
  INV_X1 U547 ( .A(n540), .ZN(n562) );
  OR2_X1 U548 ( .A1(n562), .A2(n578), .ZN(n494) );
  NOR2_X1 U549 ( .A1(n485), .A2(n494), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n491), .A2(n574), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U552 ( .A(G57GAT), .B(n488), .Z(G1332GAT) );
  NAND2_X1 U553 ( .A1(n548), .A2(n491), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n489), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U555 ( .A1(n491), .A2(n556), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n490), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U557 ( .A(G78GAT), .B(KEYINPUT43), .Z(n493) );
  NAND2_X1 U558 ( .A1(n491), .A2(n501), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n493), .B(n492), .ZN(G1335GAT) );
  NOR2_X1 U560 ( .A1(n495), .A2(n494), .ZN(n502) );
  NAND2_X1 U561 ( .A1(n574), .A2(n502), .ZN(n496) );
  XNOR2_X1 U562 ( .A(G85GAT), .B(n496), .ZN(G1336GAT) );
  XOR2_X1 U563 ( .A(G92GAT), .B(KEYINPUT109), .Z(n498) );
  NAND2_X1 U564 ( .A1(n502), .A2(n548), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(G1337GAT) );
  NAND2_X1 U566 ( .A1(n502), .A2(n556), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(KEYINPUT110), .ZN(n500) );
  XNOR2_X1 U568 ( .A(G99GAT), .B(n500), .ZN(G1338GAT) );
  NAND2_X1 U569 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(KEYINPUT44), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G106GAT), .B(n504), .ZN(G1339GAT) );
  INV_X1 U572 ( .A(n566), .ZN(n586) );
  NOR2_X1 U573 ( .A1(n546), .A2(n586), .ZN(n507) );
  NAND2_X1 U574 ( .A1(n578), .A2(n540), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n505), .B(KEYINPUT46), .ZN(n506) );
  XNOR2_X1 U576 ( .A(KEYINPUT111), .B(n508), .ZN(n510) );
  INV_X1 U577 ( .A(KEYINPUT47), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n515) );
  NOR2_X1 U579 ( .A1(n566), .A2(n589), .ZN(n511) );
  XOR2_X1 U580 ( .A(KEYINPUT45), .B(n511), .Z(n512) );
  NOR2_X1 U581 ( .A1(n581), .A2(n512), .ZN(n513) );
  NAND2_X1 U582 ( .A1(n513), .A2(n558), .ZN(n514) );
  NAND2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n516) );
  INV_X1 U584 ( .A(n549), .ZN(n518) );
  NOR2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n556), .A2(n534), .ZN(n519) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n519), .Z(n521) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U589 ( .A1(n558), .A2(n529), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  NOR2_X1 U592 ( .A1(n562), .A2(n529), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n566), .A2(n529), .ZN(n527) );
  XNOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n526) );
  XNOR2_X1 U597 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U598 ( .A(G127GAT), .B(n528), .Z(G1342GAT) );
  NOR2_X1 U599 ( .A1(n529), .A2(n570), .ZN(n533) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n531) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U602 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n577), .A2(n534), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n535), .B(KEYINPUT117), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n545), .A2(n578), .ZN(n536) );
  XNOR2_X1 U607 ( .A(n536), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n538) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n537) );
  XNOR2_X1 U610 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(n539), .Z(n542) );
  NAND2_X1 U612 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U613 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n586), .A2(n545), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n543), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n561) );
  XOR2_X1 U620 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n551) );
  NAND2_X1 U621 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U622 ( .A(n551), .B(n550), .ZN(n575) );
  INV_X1 U623 ( .A(n552), .ZN(n553) );
  OR2_X1 U624 ( .A1(n574), .A2(n553), .ZN(n554) );
  XNOR2_X1 U625 ( .A(n555), .B(KEYINPUT55), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n569) );
  NOR2_X1 U627 ( .A1(n569), .A2(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT123), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  NOR2_X1 U630 ( .A1(n562), .A2(n569), .ZN(n564) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n566), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(n567), .Z(n568) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n297), .ZN(G1351GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n573) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n580) );
  NOR2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n588) );
  INV_X1 U644 ( .A(n588), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n585), .A2(n578), .ZN(n579) );
  XOR2_X1 U646 ( .A(n580), .B(n579), .Z(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U648 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

