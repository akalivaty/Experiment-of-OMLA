//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  XOR2_X1   g000(.A(KEYINPUT24), .B(G110), .Z(new_n187));
  XNOR2_X1  g001(.A(G119), .B(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT73), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(KEYINPUT73), .ZN(new_n207));
  OAI221_X1 g021(.A(new_n189), .B1(new_n196), .B2(new_n197), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n204), .A2(G110), .B1(new_n187), .B2(new_n188), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n191), .A2(new_n193), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT74), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n211), .A2(new_n215), .A3(G146), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n209), .B(new_n210), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n219), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(KEYINPUT75), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(new_n224), .C1(new_n218), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(KEYINPUT76), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G217), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(G234), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G902), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n228), .B2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n231), .B1(new_n235), .B2(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n199), .A2(G116), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G113), .ZN(new_n246));
  INV_X1    g060(.A(G113), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT2), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT68), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n199), .A2(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(KEYINPUT2), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n245), .A2(G113), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n244), .A2(new_n249), .A3(new_n252), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n251), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n246), .B2(new_n248), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n213), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n213), .A2(G143), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT65), .B1(new_n213), .B2(G143), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n270), .B2(G146), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n213), .A2(KEYINPUT64), .A3(G143), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n201), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n272), .A2(new_n274), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n272), .A4(new_n277), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n267), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(G137), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT11), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n285), .B2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(G137), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(G131), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n201), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n263), .B2(new_n264), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n281), .A2(new_n272), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n291), .A2(G131), .ZN(new_n301));
  INV_X1    g115(.A(new_n290), .ZN(new_n302));
  OAI21_X1  g116(.A(G131), .B1(new_n302), .B2(new_n286), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n284), .A2(new_n305), .A3(new_n292), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n292), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT67), .B1(new_n284), .B2(new_n292), .ZN(new_n309));
  INV_X1    g123(.A(new_n304), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n261), .B(new_n307), .C1(new_n311), .C2(KEYINPUT30), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n284), .A2(new_n305), .A3(new_n292), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n305), .B1(new_n284), .B2(new_n292), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n310), .A2(new_n261), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT26), .B(G101), .Z(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G210), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT31), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n293), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n292), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n304), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n261), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(new_n317), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT28), .B1(new_n316), .B2(new_n293), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n323), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n312), .A2(new_n336), .A3(new_n317), .A4(new_n324), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G472), .A2(G902), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n294), .A2(new_n304), .A3(new_n306), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(new_n261), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n315), .A2(new_n316), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT28), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n349));
  INV_X1    g163(.A(new_n334), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n261), .A2(new_n345), .B1(new_n315), .B2(new_n316), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n350), .B(new_n351), .C1(new_n353), .C2(new_n327), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT72), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n355), .A3(new_n230), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n312), .A2(new_n317), .A3(new_n323), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G472), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n239), .B1(new_n344), .B2(new_n360), .ZN(new_n361));
  OAI22_X1  g175(.A1(new_n214), .A2(new_n216), .B1(new_n213), .B2(new_n212), .ZN(new_n362));
  AOI21_X1  g176(.A(G143), .B1(new_n319), .B2(G214), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT18), .A2(G131), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT18), .B(G131), .C1(new_n368), .C2(new_n363), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n196), .A2(new_n197), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT17), .B(G131), .C1(new_n368), .C2(new_n363), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT86), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n194), .A2(new_n195), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n213), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n375), .A2(new_n372), .A3(KEYINPUT86), .A4(new_n210), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n364), .A2(new_n377), .A3(new_n365), .ZN(new_n378));
  OAI21_X1  g192(.A(G131), .B1(new_n368), .B2(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n370), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n370), .B(KEYINPUT88), .C1(new_n373), .C2(new_n382), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n370), .B(new_n390), .C1(new_n373), .C2(new_n382), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n383), .B2(new_n384), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n386), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n230), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G475), .ZN(new_n398));
  NAND2_X1  g212(.A1(G234), .A2(G237), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G952), .A3(new_n220), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT21), .B(G898), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT93), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n399), .A2(G902), .A3(G953), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n270), .A2(G128), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n201), .A2(G143), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n285), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G122), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G116), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n241), .A2(G122), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G107), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G122), .ZN(new_n423));
  INV_X1    g237(.A(G107), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n417), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n201), .B2(G143), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n415), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n414), .A2(new_n427), .ZN(new_n430));
  OAI21_X1  g244(.A(G134), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n414), .A2(new_n415), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G134), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n416), .B1(new_n424), .B2(new_n423), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n241), .A2(KEYINPUT14), .A3(G122), .ZN(new_n435));
  OAI211_X1 g249(.A(G107), .B(new_n435), .C1(new_n421), .C2(KEYINPUT14), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n426), .A2(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n438), .A2(new_n229), .A3(G953), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT91), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n422), .A2(new_n425), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n431), .A3(new_n416), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n433), .A2(new_n416), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n425), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n445), .B2(new_n447), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n442), .A2(new_n444), .A3(KEYINPUT90), .A4(new_n439), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n230), .B(new_n413), .C1(new_n449), .C2(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n440), .A2(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n412), .B1(new_n455), .B2(G902), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n362), .A2(new_n367), .A3(new_n369), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n212), .A2(KEYINPUT19), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT19), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n213), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n378), .A2(new_n379), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n462), .A2(new_n210), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n391), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n393), .ZN(new_n466));
  NOR2_X1   g280(.A1(G475), .A2(G902), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT87), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n458), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AOI211_X1 g284(.A(KEYINPUT20), .B(new_n468), .C1(new_n465), .C2(new_n393), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n398), .A2(new_n407), .A3(new_n457), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n397), .B2(G475), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(KEYINPUT94), .A3(new_n407), .A4(new_n457), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G214), .B1(G237), .B2(G902), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  MUX2_X1   g295(.A(new_n300), .B(new_n284), .S(G125), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n220), .A2(G224), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n482), .A2(KEYINPUT7), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(KEYINPUT7), .B2(new_n483), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G122), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT8), .Z(new_n487));
  OAI21_X1  g301(.A(KEYINPUT79), .B1(new_n389), .B2(G107), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n424), .A3(G104), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n389), .A2(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(G101), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n424), .A3(G104), .ZN(new_n497));
  INV_X1    g311(.A(G101), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n491), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n493), .B1(new_n492), .B2(G101), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n244), .B2(new_n252), .ZN(new_n504));
  OAI21_X1  g318(.A(G113), .B1(new_n250), .B2(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n260), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n505), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n508), .A2(KEYINPUT85), .B1(new_n503), .B2(new_n258), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n260), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g326(.A(new_n487), .B(new_n507), .C1(new_n502), .C2(new_n512), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n484), .A2(new_n485), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n495), .A2(new_n497), .A3(new_n491), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT78), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n495), .A2(new_n497), .A3(new_n517), .A4(new_n491), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(G101), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n516), .A2(new_n522), .A3(G101), .A4(new_n518), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n261), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n492), .A2(G101), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT80), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n499), .A3(new_n494), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n527), .A2(new_n506), .A3(KEYINPUT82), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT82), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n258), .B1(new_n253), .B2(new_n254), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT69), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT69), .B1(new_n250), .B2(new_n251), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT5), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n533), .B2(new_n508), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n502), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n486), .B(new_n524), .C1(new_n528), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT82), .B1(new_n527), .B2(new_n506), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n494), .A2(new_n499), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n540), .A3(new_n529), .A4(new_n526), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n261), .A2(new_n523), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n539), .A2(new_n541), .B1(new_n542), .B2(new_n521), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT83), .A3(new_n486), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n486), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT6), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n537), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT83), .B1(new_n543), .B2(new_n486), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT6), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n543), .A2(new_n486), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n483), .B(KEYINPUT84), .Z(new_n555));
  XNOR2_X1  g369(.A(new_n482), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n546), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n538), .B2(new_n544), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n562), .B2(new_n547), .ZN(new_n563));
  INV_X1    g377(.A(new_n556), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n558), .A3(new_n546), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n481), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n479), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n230), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G140), .ZN(new_n573));
  INV_X1    g387(.A(G227), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(G953), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n268), .A2(new_n271), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n296), .B1(new_n578), .B2(new_n280), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(new_n299), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n580), .B2(new_n527), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n279), .A2(new_n283), .ZN(new_n582));
  INV_X1    g396(.A(new_n267), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n521), .A2(new_n582), .A3(new_n583), .A4(new_n523), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n291), .B(new_n377), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n540), .A2(new_n300), .A3(KEYINPUT10), .A4(new_n526), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n581), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n299), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n540), .A2(new_n588), .A3(new_n526), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n297), .B(new_n299), .C1(new_n500), .C2(new_n501), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT12), .B1(new_n591), .B2(new_n292), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n593), .B(new_n585), .C1(new_n589), .C2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n576), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n584), .A3(new_n586), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n292), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n576), .A2(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n572), .B1(new_n600), .B2(G469), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n592), .A2(new_n594), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n587), .A2(new_n596), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n596), .B1(new_n599), .B2(new_n587), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n571), .B(new_n230), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI211_X1 g420(.A(KEYINPUT81), .B(new_n570), .C1(new_n601), .C2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT81), .ZN(new_n608));
  INV_X1    g422(.A(new_n572), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n595), .A2(new_n576), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n597), .A2(new_n599), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(G469), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n613), .B2(new_n569), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n361), .A2(new_n568), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT95), .B(G101), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  NAND4_X1  g432(.A1(new_n565), .A2(KEYINPUT96), .A3(new_n558), .A4(new_n546), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n480), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n560), .A2(new_n621), .A3(new_n566), .ZN(new_n622));
  OR3_X1    g436(.A1(new_n437), .A2(KEYINPUT98), .A3(new_n439), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n437), .B1(KEYINPUT98), .B2(new_n439), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(KEYINPUT33), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n408), .A2(G902), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n455), .A2(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n455), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n625), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n408), .B1(new_n455), .B2(G902), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n398), .A2(new_n473), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n620), .A2(new_n622), .A3(new_n407), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n338), .A2(new_n230), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n638), .A2(G472), .B1(new_n338), .B2(new_n339), .ZN(new_n639));
  INV_X1    g453(.A(new_n239), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n615), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AOI211_X1 g458(.A(new_n472), .B(new_n457), .C1(new_n397), .C2(G475), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n620), .A2(new_n622), .A3(new_n407), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n641), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n225), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(KEYINPUT36), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(new_n218), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n232), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n237), .B2(new_n238), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n615), .A2(new_n639), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n568), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AND3_X1   g473(.A1(new_n615), .A2(new_n622), .A3(new_n620), .ZN(new_n660));
  INV_X1    g474(.A(new_n655), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n344), .B2(new_n360), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n401), .B1(new_n405), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n645), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n660), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XOR2_X1   g483(.A(new_n664), .B(KEYINPUT39), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n615), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n560), .A2(new_n566), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n673), .B(new_n674), .Z(new_n675));
  NOR4_X1   g489(.A1(new_n655), .A2(new_n457), .A3(new_n477), .A4(new_n481), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n312), .A2(new_n317), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n323), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n353), .A2(new_n323), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n230), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n342), .B1(new_n338), .B2(new_n339), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n672), .A2(new_n675), .A3(new_n676), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  NAND2_X1  g500(.A1(new_n635), .A2(new_n665), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n660), .A2(new_n662), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  OAI21_X1  g504(.A(new_n360), .B1(new_n682), .B2(new_n683), .ZN(new_n691));
  INV_X1    g505(.A(new_n604), .ZN(new_n692));
  INV_X1    g506(.A(new_n605), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n571), .B1(new_n694), .B2(new_n230), .ZN(new_n695));
  INV_X1    g509(.A(new_n606), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n570), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n640), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n637), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT101), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n647), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND3_X1   g519(.A1(new_n620), .A2(new_n622), .A3(new_n697), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n662), .A2(new_n706), .A3(new_n479), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NAND2_X1  g522(.A1(new_n638), .A2(G472), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n638), .A2(KEYINPUT102), .A3(G472), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n348), .A2(new_n350), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n326), .B(new_n337), .C1(new_n713), .C2(new_n324), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n711), .A2(new_n712), .B1(new_n339), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  INV_X1    g530(.A(new_n457), .ZN(new_n717));
  INV_X1    g531(.A(G475), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n395), .A2(new_n387), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT89), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n392), .A3(new_n393), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n721), .B2(new_n230), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n716), .B(new_n717), .C1(new_n722), .C2(new_n472), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT103), .B1(new_n477), .B2(new_n457), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(new_n724), .A3(new_n407), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n715), .A2(new_n706), .A3(new_n640), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND2_X1  g541(.A1(new_n714), .A2(new_n339), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT102), .B1(new_n638), .B2(G472), .ZN(new_n729));
  INV_X1    g543(.A(G472), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n710), .B(new_n730), .C1(new_n338), .C2(new_n230), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n655), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n620), .A2(new_n622), .A3(new_n697), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n733), .A3(new_n687), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n192), .ZN(G27));
  AOI21_X1  g549(.A(new_n570), .B1(new_n601), .B2(new_n606), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n560), .A2(new_n480), .A3(new_n566), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n361), .B(new_n688), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n737), .B(KEYINPUT104), .ZN(new_n744));
  INV_X1    g558(.A(new_n742), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n361), .A3(new_n688), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  OAI211_X1 g562(.A(new_n361), .B(new_n667), .C1(new_n738), .C2(new_n739), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n744), .A2(new_n751), .A3(new_n361), .A4(new_n667), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  NAND2_X1  g568(.A1(new_n631), .A2(new_n634), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n477), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  INV_X1    g571(.A(new_n639), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n655), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n600), .A2(KEYINPUT45), .ZN(new_n763));
  OAI21_X1  g577(.A(G469), .B1(new_n600), .B2(KEYINPUT45), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n765), .B2(new_n609), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n696), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n609), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n570), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n670), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n560), .A2(new_n480), .A3(new_n566), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT107), .Z(new_n772));
  NAND4_X1  g586(.A1(new_n761), .A2(new_n762), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  XNOR2_X1  g588(.A(new_n769), .B(KEYINPUT47), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n691), .A2(new_n771), .A3(new_n640), .A4(new_n687), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT109), .Z(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n190), .ZN(G42));
  NOR2_X1   g595(.A1(new_n695), .A2(new_n696), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n239), .A2(new_n481), .A3(new_n570), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n675), .A2(new_n787), .A3(new_n684), .A4(new_n756), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n757), .A2(new_n401), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n711), .A2(new_n712), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n640), .A3(new_n728), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n697), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n675), .A2(new_n480), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(KEYINPUT50), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n794), .A3(new_n797), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n771), .A2(new_n796), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n732), .ZN(new_n805));
  INV_X1    g619(.A(new_n684), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n803), .A3(new_n401), .A4(new_n640), .ZN(new_n807));
  INV_X1    g621(.A(new_n477), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n755), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n795), .A2(new_n772), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n775), .B1(new_n570), .B2(new_n782), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n811), .B2(KEYINPUT115), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT51), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n813), .B2(new_n814), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n691), .A2(new_n640), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n804), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT48), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n795), .A2(new_n706), .ZN(new_n824));
  INV_X1    g638(.A(G952), .ZN(new_n825));
  INV_X1    g639(.A(new_n807), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n825), .B(G953), .C1(new_n826), .C2(new_n635), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n817), .A2(new_n828), .A3(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n715), .A2(new_n706), .A3(new_n655), .A4(new_n688), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n620), .A2(new_n622), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n723), .A2(new_n724), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n654), .B(new_n665), .C1(new_n237), .C2(new_n238), .ZN(new_n836));
  INV_X1    g650(.A(new_n736), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n684), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n833), .A2(new_n668), .A3(new_n689), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT52), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n565), .A2(new_n558), .A3(new_n546), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n558), .B1(new_n565), .B2(new_n546), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n480), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n407), .B1(new_n635), .B2(new_n645), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n640), .A3(new_n615), .A4(new_n639), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n477), .A2(new_n457), .A3(new_n665), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n607), .A2(new_n614), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n771), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n691), .A2(new_n849), .A3(new_n850), .A4(new_n655), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n616), .A2(new_n657), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n715), .A2(new_n655), .A3(new_n688), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n738), .A2(new_n739), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n725), .A2(new_n622), .A3(new_n620), .A4(new_n697), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n691), .A2(new_n479), .A3(new_n655), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n793), .A2(new_n857), .B1(new_n733), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n698), .B1(new_n636), .B2(new_n646), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n856), .A2(new_n747), .A3(new_n753), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n841), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n691), .A2(new_n655), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n615), .A2(new_n620), .A3(new_n622), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(new_n666), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT111), .B1(new_n734), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n867), .A2(new_n868), .A3(new_n687), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n684), .A2(new_n838), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n835), .A2(new_n622), .A3(new_n620), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n833), .A2(new_n668), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n840), .A2(new_n875), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n700), .A2(new_n704), .A3(new_n707), .A4(new_n726), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n855), .A3(new_n852), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n746), .A2(new_n743), .B1(new_n750), .B2(new_n752), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT112), .B1(new_n885), .B2(new_n863), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n866), .B1(new_n886), .B2(new_n864), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT113), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n863), .B1(new_n841), .B2(new_n862), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(KEYINPUT53), .A3(new_n883), .A4(new_n884), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n888), .B1(new_n887), .B2(KEYINPUT54), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n831), .A2(new_n832), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n789), .B1(new_n896), .B2(new_n897), .ZN(G75));
  AOI21_X1  g712(.A(new_n230), .B1(new_n890), .B2(new_n891), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(G210), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n554), .A2(new_n556), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(new_n565), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n825), .A2(G953), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n903), .B2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(G51));
  INV_X1    g726(.A(new_n909), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n230), .B(new_n765), .C1(new_n890), .C2(new_n891), .ZN(new_n914));
  INV_X1    g728(.A(new_n694), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n892), .B2(KEYINPUT54), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n893), .B(new_n917), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n572), .B(KEYINPUT57), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n920), .B2(KEYINPUT120), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n893), .B(new_n917), .ZN(new_n922));
  INV_X1    g736(.A(new_n919), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n694), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n913), .B1(new_n921), .B2(new_n926), .ZN(G54));
  AND3_X1   g741(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n928), .B2(new_n466), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n913), .B1(new_n928), .B2(new_n466), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n928), .A2(KEYINPUT121), .A3(new_n466), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G60));
  OAI21_X1  g747(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NOR3_X1   g750(.A1(new_n922), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n936), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n894), .B2(new_n895), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n913), .B(new_n937), .C1(new_n934), .C2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n892), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n228), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n890), .B2(new_n891), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n653), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT122), .B1(new_n946), .B2(new_n909), .ZN(new_n952));
  OAI211_X1 g766(.A(KEYINPUT122), .B(new_n909), .C1(new_n947), .C2(new_n228), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n948), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n228), .B1(new_n892), .B2(new_n943), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n913), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n953), .A3(new_n948), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n960), .B2(new_n951), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n949), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n949), .C1(new_n956), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(G66));
  AOI21_X1  g780(.A(new_n220), .B1(new_n403), .B2(G224), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  AOI22_X1  g782(.A1(new_n568), .A2(new_n656), .B1(new_n641), .B2(new_n846), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n861), .A2(new_n616), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n968), .B1(new_n971), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n554), .B1(G898), .B2(new_n220), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  OAI21_X1  g788(.A(new_n307), .B1(new_n311), .B2(KEYINPUT30), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n460), .A2(new_n461), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n870), .A2(new_n689), .A3(new_n878), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n685), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g794(.A(new_n671), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n850), .C1(new_n635), .C2(new_n645), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n773), .B1(new_n820), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n780), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(KEYINPUT62), .B2(new_n979), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n977), .B1(new_n985), .B2(new_n220), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n780), .B1(new_n752), .B2(new_n750), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n770), .A2(new_n361), .A3(new_n834), .A4(new_n835), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n773), .A2(new_n747), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n987), .A2(new_n220), .A3(new_n978), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(G900), .A2(G953), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n977), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n986), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(G953), .B1(new_n574), .B2(new_n663), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G72));
  NAND4_X1  g809(.A1(new_n987), .A2(new_n971), .A3(new_n978), .A4(new_n989), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n358), .B(KEYINPUT126), .Z(new_n1000));
  AOI21_X1  g814(.A(new_n913), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n887), .ZN(new_n1002));
  INV_X1    g816(.A(new_n678), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n358), .A3(new_n998), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n998), .B1(new_n985), .B2(new_n970), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n678), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1001), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT127), .ZN(G57));
endmodule


