//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n198), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT0), .B(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n207), .B(new_n212), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G104), .B(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT73), .B1(new_n215), .B2(new_n195), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n193), .A2(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n196), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G101), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n216), .A2(new_n220), .B1(new_n221), .B2(new_n195), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n223), .A2(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n226), .A2(new_n203), .A3(new_n205), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n201), .A2(new_n214), .B1(new_n222), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  INV_X1    g046(.A(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G137), .ZN(new_n234));
  INV_X1    g048(.A(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT11), .A3(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n234), .A2(new_n236), .A3(new_n240), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n203), .A2(new_n205), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(KEYINPUT1), .C1(new_n204), .C2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n208), .A2(new_n226), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n222), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT75), .B1(new_n252), .B2(new_n229), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n254));
  AOI211_X1 g068(.A(new_n254), .B(KEYINPUT10), .C1(new_n222), .C2(new_n251), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n231), .B(new_n243), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n219), .B1(new_n218), .B2(G101), .ZN(new_n257));
  AOI211_X1 g071(.A(KEYINPUT73), .B(new_n195), .C1(new_n217), .C2(new_n196), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n197), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n223), .A2(KEYINPUT74), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G128), .A3(new_n246), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n227), .B1(new_n261), .B2(new_n244), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n223), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n244), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n250), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n222), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n242), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n242), .A2(KEYINPUT76), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(KEYINPUT12), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(KEYINPUT12), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(new_n242), .C1(new_n263), .C2(new_n267), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n256), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G140), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n231), .B1(new_n253), .B2(new_n255), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n242), .ZN(new_n280));
  INV_X1    g094(.A(new_n277), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n256), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(G469), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G469), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n289));
  INV_X1    g103(.A(new_n256), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n254), .B1(new_n263), .B2(KEYINPUT10), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n252), .A2(KEYINPUT75), .A3(new_n229), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n243), .B1(new_n293), .B2(new_n231), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n256), .A2(new_n270), .A3(new_n281), .A4(new_n272), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n288), .A2(new_n289), .B1(new_n297), .B2(new_n284), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n284), .B1(new_n273), .B2(new_n277), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n289), .B(new_n286), .C1(new_n299), .C2(new_n282), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n213), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  OR2_X1    g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n204), .A2(G146), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n202), .A2(G143), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n212), .B1(new_n308), .B2(new_n207), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n242), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n233), .A2(G137), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n235), .A2(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n266), .A2(new_n241), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G113), .ZN(new_n317));
  INV_X1    g131(.A(G113), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT65), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G116), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(G113), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n320), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n327), .ZN(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n241), .A2(new_n313), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n228), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n210), .B1(new_n241), .B2(new_n239), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n315), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n332), .B1(KEYINPUT65), .B2(new_n331), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT2), .B(G113), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT66), .B1(new_n325), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n329), .A2(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n310), .A2(new_n314), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n350));
  INV_X1    g164(.A(G210), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n351), .A2(G237), .A3(G953), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G101), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n315), .A2(new_n357), .A3(new_n336), .A4(new_n341), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n343), .A2(new_n349), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT31), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n358), .A2(new_n349), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT31), .A3(new_n356), .A4(new_n343), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n211), .A2(new_n213), .B1(new_n241), .B2(new_n239), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n365), .A2(new_n339), .A3(new_n336), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n242), .A2(new_n207), .A3(new_n308), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n348), .B1(new_n367), .B2(new_n314), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n355), .B(KEYINPUT70), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n349), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT71), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n314), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n336), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n376), .B2(new_n349), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n369), .B(new_n370), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n364), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(G472), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT32), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT32), .ZN(new_n382));
  INV_X1    g196(.A(new_n378), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n361), .B2(new_n363), .ZN(new_n384));
  INV_X1    g198(.A(new_n380), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n369), .B1(new_n374), .B2(new_n377), .ZN(new_n387));
  INV_X1    g201(.A(new_n370), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n358), .A2(new_n349), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n355), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n348), .B1(new_n310), .B2(new_n314), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n366), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n372), .B1(new_n396), .B2(new_n371), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n355), .A2(new_n393), .ZN(new_n399));
  AOI21_X1  g213(.A(G902), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G472), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n381), .A2(new_n386), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n321), .B2(G128), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n405), .B(new_n406), .C1(G119), .C2(new_n225), .ZN(new_n407));
  XNOR2_X1  g221(.A(G119), .B(G128), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT24), .B(G110), .Z(new_n409));
  AOI22_X1  g223(.A1(new_n407), .A2(G110), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G125), .B(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT16), .ZN(new_n413));
  INV_X1    g227(.A(G140), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G125), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(G146), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G146), .B1(new_n412), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n407), .A2(G110), .B1(new_n408), .B2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n411), .A2(new_n202), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT22), .B(G137), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(new_n422), .A3(new_n426), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT25), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n285), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n285), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT25), .ZN(new_n434));
  NAND2_X1  g248(.A1(G217), .A2(G902), .ZN(new_n435));
  INV_X1    g249(.A(G217), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(G234), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G237), .A2(G953), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n444), .A2(G143), .A3(G214), .ZN(new_n445));
  AOI21_X1  g259(.A(G143), .B1(new_n444), .B2(G214), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT18), .A2(G131), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n414), .A2(G125), .ZN(new_n451));
  INV_X1    g265(.A(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G146), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n421), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n445), .A2(new_n446), .A3(G131), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(G214), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n204), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n444), .A2(G143), .A3(G214), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n240), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n458), .A2(new_n462), .A3(KEYINPUT17), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n415), .B1(new_n454), .B2(new_n413), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n202), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n445), .B2(new_n446), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n465), .B(new_n416), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G113), .B(G122), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n190), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n457), .B(new_n471), .C1(new_n463), .C2(new_n468), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n285), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G475), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n458), .B2(new_n462), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n460), .A2(new_n240), .A3(new_n461), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n467), .A2(new_n481), .A3(KEYINPUT84), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n411), .A2(KEYINPUT19), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n411), .A2(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n202), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n416), .A3(new_n482), .A4(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(new_n457), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n474), .B1(new_n487), .B2(new_n471), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n471), .B1(new_n486), .B2(new_n457), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n478), .B(new_n489), .C1(new_n475), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n477), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n496));
  OAI21_X1  g310(.A(G134), .B1(new_n496), .B2(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n225), .A2(G143), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n496), .A2(KEYINPUT85), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n225), .B2(G143), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n204), .A2(G128), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n498), .A3(new_n233), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G116), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n323), .A2(G122), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(new_n507), .A3(new_n193), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n193), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n495), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n503), .A2(new_n498), .A3(new_n233), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n507), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G107), .ZN(new_n514));
  XNOR2_X1  g328(.A(G116), .B(G122), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n193), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n501), .A2(new_n496), .A3(KEYINPUT85), .A4(new_n498), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(G134), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(KEYINPUT86), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n233), .B1(new_n503), .B2(new_n498), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n516), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n323), .A2(KEYINPUT14), .A3(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n515), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n523), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n503), .A2(new_n498), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G134), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n504), .ZN(new_n533));
  OAI211_X1 g347(.A(G107), .B(new_n526), .C1(new_n513), .C2(KEYINPUT14), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT87), .A4(new_n516), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n187), .A2(new_n436), .A3(G953), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n522), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n522), .B2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n285), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(G478), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n522), .A2(new_n536), .ZN(new_n544));
  INV_X1    g358(.A(new_n537), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n538), .ZN(new_n547));
  INV_X1    g361(.A(G478), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(new_n285), .C1(KEYINPUT15), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(G234), .A2(G237), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(G952), .A3(new_n275), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n550), .A2(G902), .A3(G953), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT21), .B(G898), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT88), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n543), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n494), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n323), .A2(G119), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT5), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n318), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n334), .B2(new_n335), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT78), .B1(new_n565), .B2(new_n259), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n198), .A2(G101), .A3(new_n199), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n336), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n346), .A2(new_n347), .B1(new_n560), .B2(new_n563), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n222), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G122), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT79), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n579), .A3(new_n574), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n576), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n566), .A2(new_n569), .A3(new_n572), .A4(new_n575), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT80), .B1(new_n266), .B2(G125), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n210), .A2(G125), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n228), .A2(new_n587), .A3(new_n452), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G224), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G953), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n584), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G210), .B1(G237), .B2(G902), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT7), .B1(new_n590), .B2(G953), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT82), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n589), .A2(new_n595), .ZN(new_n599));
  OAI21_X1  g413(.A(G113), .B1(new_n322), .B2(KEYINPUT5), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n601), .A2(new_n560), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n334), .A2(new_n335), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n222), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n575), .B(KEYINPUT8), .Z(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n570), .B2(new_n259), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n599), .A2(new_n583), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n598), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n593), .A2(new_n594), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n594), .B(KEYINPUT83), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n593), .B2(new_n610), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n558), .B(new_n559), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n302), .A2(new_n403), .A3(new_n443), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(G472), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n379), .B2(new_n285), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n384), .A2(G902), .A3(new_n620), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n302), .A2(new_n443), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n539), .B2(new_n540), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n548), .A2(G902), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT91), .B1(new_n544), .B2(new_n545), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n630), .B(new_n537), .C1(new_n522), .C2(new_n536), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT92), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n538), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n522), .A2(new_n536), .A3(KEYINPUT92), .A4(new_n537), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(KEYINPUT33), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n627), .B(new_n628), .C1(new_n632), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n541), .A2(new_n548), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n637), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT93), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n494), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(KEYINPUT94), .B(new_n494), .C1(new_n639), .C2(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n593), .A2(new_n610), .ZN(new_n647));
  INV_X1    g461(.A(new_n594), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT90), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n593), .A2(new_n594), .A3(new_n610), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n593), .A2(KEYINPUT90), .A3(new_n594), .A4(new_n610), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n559), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n654), .A3(new_n556), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n625), .A2(new_n646), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT34), .B(G104), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  AOI21_X1  g472(.A(new_n494), .B1(new_n543), .B2(new_n549), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n556), .A2(new_n652), .A3(new_n654), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n625), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n423), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n440), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n439), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n615), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n302), .A3(new_n624), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AOI21_X1  g488(.A(new_n385), .B1(new_n364), .B2(new_n378), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n675), .A2(KEYINPUT32), .B1(new_n401), .B2(G472), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n670), .B1(new_n676), .B2(new_n386), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n543), .A2(new_n549), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n552), .B1(new_n553), .B2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n494), .A3(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n652), .A2(new_n654), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n682), .A3(new_n302), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n685));
  INV_X1    g499(.A(new_n296), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n281), .B1(new_n280), .B2(new_n256), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n284), .B(new_n285), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n286), .B1(new_n299), .B2(new_n282), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(KEYINPUT77), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n188), .B1(new_n690), .B2(new_n300), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n680), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n685), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n298), .A2(new_n301), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(KEYINPUT40), .A3(new_n188), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT97), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n694), .A2(new_n696), .A3(KEYINPUT97), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n647), .A2(new_n612), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n651), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n702), .B(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n359), .B1(new_n388), .B2(new_n396), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n285), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G472), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n381), .A2(new_n386), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n543), .A2(new_n549), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n494), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n668), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n559), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n705), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n699), .A2(new_n700), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT98), .B(G143), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G45));
  NAND2_X1  g532(.A1(new_n651), .A2(new_n650), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n594), .B1(new_n593), .B2(new_n610), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n559), .B(new_n653), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n680), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n494), .B(new_n722), .C1(new_n639), .C2(new_n640), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n677), .A2(new_n724), .A3(new_n302), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT99), .B(G146), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G48));
  AOI21_X1  g541(.A(new_n442), .B1(new_n676), .B2(new_n386), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n652), .A2(new_n556), .A3(new_n654), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n285), .B1(new_n686), .B2(new_n687), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n188), .A3(new_n688), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n728), .A2(new_n645), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT41), .B(G113), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n734), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n660), .A2(new_n728), .A3(new_n733), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  INV_X1    g553(.A(new_n558), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n721), .A2(new_n740), .A3(new_n732), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n677), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  OAI21_X1  g557(.A(G472), .B1(new_n384), .B2(G902), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n397), .A2(new_n370), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n364), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n380), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n747), .A3(new_n443), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n744), .A2(new_n747), .A3(KEYINPUT101), .A4(new_n443), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n731), .A2(new_n188), .A3(new_n688), .A4(new_n556), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n494), .A2(new_n711), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n721), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  NAND3_X1  g571(.A1(new_n744), .A2(new_n747), .A3(new_n668), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n723), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n721), .A2(new_n732), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  XOR2_X1   g576(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n763));
  NAND2_X1  g577(.A1(new_n688), .A2(new_n287), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n278), .A2(KEYINPUT102), .A3(new_n282), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT102), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n273), .A2(new_n766), .A3(new_n277), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n284), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n188), .B1(new_n764), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n701), .A2(new_n559), .A3(new_n651), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n728), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n763), .B1(new_n772), .B2(new_n723), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n386), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n386), .A2(new_n774), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n676), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n723), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n443), .A3(new_n771), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND3_X1  g596(.A1(new_n728), .A2(new_n771), .A3(new_n681), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NOR2_X1   g598(.A1(new_n624), .A2(new_n713), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n639), .A2(new_n640), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n786), .B(KEYINPUT43), .C1(new_n787), .C2(new_n494), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  INV_X1    g603(.A(new_n640), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n637), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n494), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n789), .B1(new_n792), .B2(KEYINPUT107), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT108), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n788), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT44), .B1(new_n796), .B2(new_n785), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n770), .ZN(new_n798));
  AOI211_X1 g612(.A(G469), .B(G902), .C1(new_n295), .C2(new_n296), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT106), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n273), .A2(new_n766), .A3(new_n277), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n766), .B1(new_n273), .B2(new_n277), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n282), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n765), .A2(new_n767), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(KEYINPUT106), .A3(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(KEYINPUT45), .A2(G469), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n283), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT105), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n287), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT46), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n799), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT106), .B1(new_n806), .B2(KEYINPUT45), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n800), .B(new_n804), .C1(new_n765), .C2(new_n767), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT105), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n810), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(KEYINPUT46), .A3(new_n287), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n189), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n795), .A2(new_n798), .A3(new_n692), .A4(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT109), .B(G137), .Z(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(G39));
  NAND2_X1  g639(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n286), .B1(new_n817), .B2(new_n819), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n688), .B1(new_n827), .B2(KEYINPUT46), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n812), .A2(new_n813), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n188), .B(new_n826), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n403), .A2(new_n723), .A3(new_n770), .A4(new_n443), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n832));
  OAI211_X1 g646(.A(new_n830), .B(new_n831), .C1(new_n822), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  AND3_X1   g648(.A1(new_n793), .A2(new_n552), .A3(new_n788), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n752), .ZN(new_n836));
  INV_X1    g650(.A(new_n770), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n830), .B1(new_n822), .B2(new_n832), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n297), .A2(new_n284), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n799), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n189), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n732), .A2(new_n770), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n710), .A2(new_n844), .A3(new_n443), .A4(new_n552), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n845), .A2(new_n494), .A3(new_n640), .A4(new_n639), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n835), .A2(new_n844), .ZN(new_n847));
  INV_X1    g661(.A(new_n758), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n732), .A2(new_n559), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n835), .A2(new_n705), .A3(new_n752), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT115), .B(new_n858), .C1(new_n843), .C2(new_n855), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n777), .A2(new_n443), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n847), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n860), .B(KEYINPUT48), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(G952), .B(new_n275), .C1(new_n845), .C2(new_n646), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n836), .B2(new_n760), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n857), .A2(new_n859), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n756), .A2(new_n734), .A3(new_n738), .A4(new_n742), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT111), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n403), .A2(new_n733), .A3(new_n443), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n752), .A2(new_n755), .B1(new_n876), .B2(new_n660), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n655), .B1(new_n643), .B2(new_n644), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n878), .A2(new_n876), .B1(new_n677), .B2(new_n741), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n683), .A2(new_n761), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n683), .A2(new_n761), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n652), .A2(new_n654), .A3(new_n712), .ZN(new_n887));
  INV_X1    g701(.A(new_n434), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n438), .B1(new_n433), .B2(KEYINPUT25), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n667), .B(new_n722), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n439), .A2(KEYINPUT114), .A3(new_n667), .A4(new_n722), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n188), .C1(new_n764), .C2(new_n768), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n887), .A2(new_n896), .A3(new_n709), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(KEYINPUT52), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n884), .A2(new_n725), .A3(new_n886), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n725), .A2(new_n683), .A3(new_n761), .A4(new_n897), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(new_n783), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n773), .B2(new_n780), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n641), .B1(new_n494), .B2(new_n678), .ZN(new_n907));
  INV_X1    g721(.A(new_n559), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n701), .B2(new_n651), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n909), .A3(new_n556), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n617), .B(new_n672), .C1(new_n625), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n759), .A2(new_n771), .ZN(new_n912));
  INV_X1    g726(.A(new_n670), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n302), .A2(new_n403), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT112), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n543), .A2(new_n549), .A3(new_n722), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n494), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n770), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n611), .A2(new_n614), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT112), .A3(new_n559), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n912), .B1(new_n914), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n911), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n906), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n882), .A2(new_n903), .A3(new_n904), .A4(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n875), .A2(new_n881), .A3(new_n906), .A4(new_n924), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n900), .B(KEYINPUT52), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT53), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n929), .A3(KEYINPUT54), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n904), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n874), .A2(new_n904), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n903), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n930), .B1(KEYINPUT54), .B2(new_n934), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n873), .A2(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n841), .B(KEYINPUT49), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n792), .A2(new_n443), .A3(new_n188), .A4(new_n559), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n939), .A3(new_n710), .A4(new_n705), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(G75));
  NAND4_X1  g755(.A1(new_n934), .A2(KEYINPUT118), .A3(G902), .A4(new_n612), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n581), .A2(new_n584), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n592), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n285), .B1(new_n931), .B2(new_n933), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT118), .B1(new_n949), .B2(new_n612), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n275), .A2(G952), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT56), .B1(new_n949), .B2(G210), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n945), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n951), .A2(new_n955), .ZN(G51));
  XNOR2_X1  g770(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n286), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT54), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n931), .A2(new_n959), .A3(new_n933), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n931), .B2(new_n933), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n295), .A2(new_n296), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n820), .B(KEYINPUT120), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n949), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n952), .B1(new_n964), .B2(new_n966), .ZN(G54));
  AND2_X1   g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n949), .A2(new_n488), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n488), .B1(new_n949), .B2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n952), .ZN(G60));
  NOR2_X1   g785(.A1(new_n632), .A2(new_n636), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n626), .B2(new_n547), .ZN(new_n973));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n973), .B(new_n975), .C1(new_n960), .C2(new_n961), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n935), .B2(new_n975), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(G63));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n435), .B(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n931), .B2(new_n933), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n666), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n953), .B1(new_n982), .B2(new_n430), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n982), .A2(new_n430), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(KEYINPUT61), .A3(new_n953), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G66));
  INV_X1    g803(.A(new_n554), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n275), .B1(new_n990), .B2(G224), .ZN(new_n991));
  INV_X1    g805(.A(new_n911), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n882), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(new_n275), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n943), .B1(G898), .B2(new_n275), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT121), .Z(new_n996));
  XNOR2_X1  g810(.A(new_n994), .B(new_n996), .ZN(G69));
  AOI21_X1  g811(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT123), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n315), .A2(new_n341), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n483), .A2(new_n484), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n677), .A2(new_n724), .A3(new_n302), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n883), .B2(KEYINPUT113), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n716), .A2(new_n1006), .A3(new_n886), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT122), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1007), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n716), .A2(new_n1006), .A3(new_n1013), .A4(new_n886), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n907), .A2(new_n837), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n728), .A3(new_n302), .A4(new_n692), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n823), .A2(new_n833), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1004), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1002), .B1(G900), .B2(new_n275), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n812), .A2(new_n813), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(new_n688), .A3(new_n821), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n777), .A2(new_n443), .A3(new_n887), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1022), .A2(new_n188), .A3(new_n692), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT124), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n822), .A2(new_n1026), .A3(new_n692), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n906), .A2(new_n886), .A3(new_n1006), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1028), .A2(new_n823), .A3(new_n833), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1020), .B1(new_n1030), .B2(new_n275), .ZN(new_n1031));
  OAI211_X1 g845(.A(KEYINPUT125), .B(new_n999), .C1(new_n1019), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n275), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1020), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1007), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1036));
  AOI21_X1  g850(.A(KEYINPUT122), .B1(new_n1007), .B2(KEYINPUT62), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1003), .B1(new_n1038), .B2(new_n1017), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1032), .A2(new_n1042), .ZN(G72));
  NOR2_X1   g857(.A1(new_n390), .A2(new_n391), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1044), .A2(new_n355), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1038), .A2(new_n993), .A3(new_n1017), .ZN(new_n1046));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1045), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1048), .B1(new_n1030), .B2(new_n993), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1051), .A2(new_n355), .A3(new_n1044), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n359), .A2(KEYINPUT126), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(new_n392), .Z(new_n1054));
  NOR2_X1   g868(.A1(new_n1054), .A2(new_n1049), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n926), .A2(new_n929), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(KEYINPUT127), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT127), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n926), .A2(new_n929), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n952), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g874(.A1(new_n1050), .A2(new_n1052), .A3(new_n1060), .ZN(G57));
endmodule


