//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT70), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n463), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2104), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n477), .A2(new_n471), .A3(KEYINPUT68), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT68), .B1(new_n477), .B2(new_n471), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n468), .A2(G2104), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n477), .A2(new_n471), .A3(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT69), .A3(G125), .ZN(new_n489));
  NAND2_X1  g064(.A1(G113), .A2(G2104), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n482), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n476), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(G160));
  NAND4_X1  g069(.A1(new_n473), .A2(new_n469), .A3(G2105), .A4(new_n471), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  XOR2_X1   g072(.A(new_n497), .B(KEYINPUT72), .Z(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G112), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n474), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G136), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G162));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n473), .A2(new_n469), .A3(new_n471), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n478), .A2(new_n479), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n505), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n463), .A2(G114), .ZN(new_n513));
  OAI21_X1  g088(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT73), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT73), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n496), .A2(G126), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  OAI21_X1  g106(.A(G543), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  INV_X1    g107(.A(G50), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n525), .A2(new_n534), .ZN(G166));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT6), .B(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .A3(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  INV_X1    g116(.A(new_n530), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(KEYINPUT75), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(G52), .B2(new_n540), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n542), .A2(G90), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n527), .A2(new_n526), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(G651), .A2(new_n560), .B1(new_n542), .B2(G81), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n540), .A2(G43), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n530), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n522), .A2(new_n538), .A3(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(G91), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT78), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n527), .A2(new_n526), .A3(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n520), .B2(new_n521), .ZN(new_n577));
  OAI21_X1  g152(.A(G65), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT9), .B1(new_n532), .B2(new_n581), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n532), .A2(KEYINPUT9), .A3(new_n581), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n580), .A2(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n574), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G166), .ZN(G303));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n524), .B1(new_n558), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n532), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(G49), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n571), .A2(G87), .A3(new_n572), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n571), .A2(G86), .A3(new_n572), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(G48), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  OAI21_X1  g170(.A(G61), .B1(new_n527), .B2(new_n526), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n595), .B1(new_n598), .B2(G651), .ZN(new_n599));
  AOI211_X1 g174(.A(KEYINPUT80), .B(new_n524), .C1(new_n596), .C2(new_n597), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n593), .B(new_n594), .C1(new_n599), .C2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n558), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(G651), .A2(new_n604), .B1(new_n542), .B2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n540), .A2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n571), .A2(G92), .A3(new_n572), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n571), .A2(KEYINPUT10), .A3(G92), .A4(new_n572), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT81), .B(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n575), .B2(new_n577), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G54), .B2(new_n540), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n613), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n608), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n608), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G286), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G299), .B(KEYINPUT83), .Z(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G297));
  AOI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G280));
  AND3_X1   g205(.A1(new_n613), .A2(new_n618), .A3(new_n621), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n621), .B1(new_n613), .B2(new_n618), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(G559), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(G148));
  NOR2_X1   g211(.A1(new_n563), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n623), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n637), .B1(new_n639), .B2(G868), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT85), .ZN(G323));
  XOR2_X1   g216(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n642));
  XNOR2_X1  g217(.A(G323), .B(new_n642), .ZN(G282));
  NAND2_X1  g218(.A1(new_n488), .A2(new_n465), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  OR2_X1    g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n651));
  INV_X1    g226(.A(G123), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n495), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n502), .B2(G135), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(KEYINPUT14), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n660), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(G401));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n647), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2096), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT19), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  INV_X1    g269(.A(new_n691), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n686), .A2(new_n687), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n688), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n694), .B(new_n698), .C1(new_n695), .C2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT99), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT26), .ZN(new_n711));
  INV_X1    g286(.A(G129), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n495), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n465), .A2(G105), .ZN(new_n714));
  INV_X1    g289(.A(G141), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n474), .B2(new_n715), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n713), .A2(KEYINPUT100), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT100), .B1(new_n713), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(KEYINPUT101), .C1(G29), .C2(G32), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT101), .B2(new_n721), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n727), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT102), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1966), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  INV_X1    g313(.A(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n463), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n495), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n502), .B2(G140), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n736), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n731), .A2(new_n735), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G35), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n748), .A2(KEYINPUT105), .A3(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(KEYINPUT105), .B1(new_n748), .B2(G29), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G162), .C2(new_n736), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT106), .B(KEYINPUT29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n727), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n623), .B2(new_n727), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G1348), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n726), .A2(new_n747), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  XOR2_X1   g334(.A(KEYINPUT103), .B(G28), .Z(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n654), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT91), .B(G16), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G19), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n563), .B2(new_n765), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n763), .B1(new_n736), .B2(new_n764), .C1(new_n767), .C2(G1341), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G1341), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n734), .A2(G1966), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n769), .B(new_n773), .C1(new_n774), .C2(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n765), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT107), .B(KEYINPUT23), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT98), .B(KEYINPUT24), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(new_n736), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n492), .B(KEYINPUT71), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n736), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n775), .B(new_n782), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n756), .A2(G1348), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n753), .A2(G2090), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n790), .B(new_n791), .C1(new_n725), .C2(new_n723), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n736), .A2(G33), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n502), .A2(G139), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n488), .A2(G127), .ZN(new_n797));
  NAND2_X1  g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n463), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n796), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n793), .B1(new_n803), .B2(new_n736), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT97), .ZN(new_n805));
  INV_X1    g380(.A(G2072), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(new_n783), .B2(new_n788), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n758), .A2(new_n789), .A3(new_n792), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n736), .A2(G25), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n502), .A2(G131), .ZN(new_n811));
  INV_X1    g386(.A(G119), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n463), .A2(G107), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n495), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n736), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n765), .A2(G24), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT92), .ZN(new_n823));
  INV_X1    g398(.A(G290), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n765), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n820), .A2(new_n821), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G23), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n830));
  NAND2_X1  g405(.A1(G288), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT93), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n829), .B1(new_n833), .B2(G16), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT33), .B(G1976), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n765), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(G22), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n837), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT94), .B(G1971), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n727), .A2(G6), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G305), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT32), .B(G1981), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n845), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n841), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT95), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n836), .A2(new_n851), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT34), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n828), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(KEYINPUT34), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT36), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n859), .A3(new_n856), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n809), .B1(new_n858), .B2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n860), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n758), .A2(new_n789), .A3(new_n792), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n808), .ZN(G150));
  NOR2_X1   g439(.A1(new_n633), .A2(new_n638), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n540), .A2(G55), .ZN(new_n867));
  NAND2_X1  g442(.A1(G80), .A2(G543), .ZN(new_n868));
  INV_X1    g443(.A(G67), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n558), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G651), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n542), .A2(G93), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n563), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n561), .A2(new_n562), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n866), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n866), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n884), .A3(new_n634), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n873), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT108), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G145));
  NAND2_X1  g467(.A1(new_n719), .A2(new_n803), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n713), .A2(new_n716), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n801), .B2(new_n802), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n518), .B(new_n743), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(new_n816), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n496), .A2(G130), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n463), .A2(G118), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n900));
  INV_X1    g475(.A(G142), .ZN(new_n901));
  OAI221_X1 g476(.A(new_n898), .B1(new_n899), .B2(new_n900), .C1(new_n901), .C2(new_n474), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n645), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n896), .A2(new_n816), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n897), .B2(new_n904), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n893), .B(new_n895), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n893), .A2(new_n895), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n787), .A2(new_n654), .ZN(new_n912));
  NAND2_X1  g487(.A1(G160), .A2(new_n764), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(G162), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(G162), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n908), .A2(new_n911), .A3(new_n914), .A4(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n917), .A2(new_n914), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n921), .A2(KEYINPUT110), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n921), .A2(KEYINPUT110), .B1(new_n911), .B2(new_n908), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT40), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT40), .B1(new_n920), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(G395));
  NAND2_X1  g502(.A1(new_n873), .A2(new_n626), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n929));
  XOR2_X1   g504(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n833), .A2(G305), .ZN(new_n932));
  XNOR2_X1  g507(.A(G303), .B(G290), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n833), .A2(G305), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n934), .ZN(new_n939));
  INV_X1    g514(.A(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n930), .A3(new_n935), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(G299), .A2(new_n619), .ZN(new_n945));
  NAND2_X1  g520(.A1(G299), .A2(new_n619), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT41), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n950), .A3(new_n946), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n639), .A2(new_n881), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n623), .A2(new_n878), .A3(new_n638), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n947), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT111), .A3(new_n950), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n953), .A3(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n929), .B1(new_n944), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n943), .A2(new_n958), .A3(KEYINPUT113), .A4(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n944), .A2(new_n960), .A3(KEYINPUT114), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT114), .B1(new_n944), .B2(new_n960), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n928), .B1(new_n966), .B2(new_n626), .ZN(G295));
  OAI21_X1  g542(.A(new_n928), .B1(new_n966), .B2(new_n626), .ZN(G331));
  NAND2_X1  g543(.A1(new_n878), .A2(G168), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n875), .A2(G286), .A3(new_n877), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(G171), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G171), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n952), .A2(new_n973), .A3(new_n957), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n941), .A2(new_n935), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n956), .B1(new_n971), .B2(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n941), .A2(KEYINPUT115), .A3(new_n935), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n974), .A2(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n951), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n973), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n948), .A2(new_n985), .A3(new_n951), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n976), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n981), .A2(new_n982), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n978), .A4(new_n977), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n984), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n979), .B2(new_n983), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(KEYINPUT43), .A3(new_n978), .A4(new_n977), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n995), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1001), .B(new_n476), .C1(new_n491), .C2(G2105), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n512), .B2(new_n517), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n488), .A2(new_n510), .B1(KEYINPUT4), .B2(new_n507), .ZN(new_n1007));
  INV_X1    g582(.A(new_n516), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT73), .ZN(new_n1009));
  INV_X1    g584(.A(G126), .ZN(new_n1010));
  OAI22_X1  g585(.A1(new_n1008), .A2(new_n1009), .B1(new_n495), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n1012), .B2(KEYINPUT117), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1002), .A2(new_n1005), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1996), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n894), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1005), .ZN(new_n1020));
  INV_X1    g595(.A(G125), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n486), .B2(new_n487), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n490), .B1(new_n1022), .B2(KEYINPUT69), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n480), .A2(new_n481), .ZN(new_n1024));
  OAI21_X1  g599(.A(G2105), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n476), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(G40), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n743), .B(G2067), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n719), .B2(G1996), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1018), .A2(new_n1019), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n816), .A2(new_n819), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n816), .A2(new_n819), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n824), .A2(new_n826), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT118), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n826), .B2(new_n824), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1028), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n518), .A2(new_n1042), .A3(new_n1006), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n492), .A2(new_n1041), .A3(new_n1043), .A4(G40), .ZN(new_n1044));
  INV_X1    g619(.A(G1956), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1012), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1002), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1052));
  OR2_X1    g627(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1046), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1348), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1044), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1002), .A2(new_n745), .A3(new_n1003), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n623), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1055), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n623), .A2(KEYINPUT124), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n623), .B2(KEYINPUT124), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n1068), .A3(new_n1058), .A4(new_n1057), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT124), .B1(new_n631), .B2(new_n632), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1057), .A2(KEYINPUT60), .A3(new_n1070), .A4(new_n1058), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n623), .A2(KEYINPUT124), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n1065), .A2(new_n1069), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1071), .A2(new_n1072), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1065), .B1(new_n1076), .B2(new_n1069), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1063), .A2(new_n1054), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT61), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1063), .A2(new_n1081), .A3(new_n1054), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1025), .A2(new_n1003), .A3(G40), .A4(new_n1026), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(KEYINPUT123), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n492), .A2(new_n1049), .A3(new_n1047), .A4(G40), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(G1996), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT123), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n563), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n563), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1080), .A2(new_n1082), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1064), .B1(new_n1078), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1027), .ZN(new_n1098));
  INV_X1    g673(.A(G2090), .ZN(new_n1099));
  INV_X1    g674(.A(G1971), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1098), .A2(new_n1099), .B1(new_n1086), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G8), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n542), .A2(G86), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n594), .B(new_n1105), .C1(new_n599), .C2(new_n600), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(G1981), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G305), .A2(G1981), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(G1981), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(G8), .A4(new_n1083), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n831), .A2(G1976), .A3(new_n832), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1083), .A2(G8), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT52), .ZN(new_n1115));
  INV_X1    g690(.A(G1976), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(G288), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1083), .A2(G8), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1112), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1086), .A2(new_n1100), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1002), .A2(new_n1099), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1096), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1103), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1966), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1086), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1002), .A2(new_n783), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1129), .B2(G286), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1098), .A2(new_n783), .B1(new_n1086), .B2(new_n1126), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G168), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT51), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1102), .B1(new_n1131), .B2(G168), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1125), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1086), .B2(G2078), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1044), .A2(new_n730), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1139), .B(G2078), .C1(new_n1003), .C2(KEYINPUT45), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1020), .A2(new_n1142), .A3(new_n1002), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1002), .A2(new_n772), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1146), .A2(new_n1139), .B1(new_n730), .B2(new_n1044), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1002), .A3(new_n1049), .ZN(new_n1148));
  AOI21_X1  g723(.A(G301), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1138), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1144), .A2(G171), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(G301), .A3(new_n1148), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT54), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1137), .B(new_n1150), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1094), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1129), .A2(G286), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1135), .B1(new_n1134), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1130), .A2(KEYINPUT51), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1133), .A2(new_n1162), .A3(new_n1136), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1149), .A2(new_n1103), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G288), .A2(G1976), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT120), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1108), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1102), .B(new_n1169), .C1(new_n1003), .C2(new_n1002), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1124), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1119), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  NAND2_X1  g748(.A1(G168), .A2(G8), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT121), .B1(new_n1129), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1177), .B(new_n1174), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1179), .A2(new_n1119), .A3(new_n1124), .A4(new_n1103), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1173), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1177), .B1(new_n1131), .B2(new_n1174), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1129), .A2(KEYINPUT121), .A3(new_n1175), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1181), .B(new_n1173), .C1(new_n1125), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1165), .B(new_n1172), .C1(new_n1182), .C2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1040), .B1(new_n1157), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1028), .A2(new_n1015), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT46), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1029), .A2(new_n894), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1028), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(KEYINPUT47), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1194), .A2(KEYINPUT47), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1035), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1037), .A2(new_n1028), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1195), .A2(new_n1196), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n743), .A2(new_n745), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT127), .B(new_n1028), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1204), .B1(new_n1205), .B2(new_n1014), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1200), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1189), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g783(.A1(new_n920), .A2(new_n924), .ZN(new_n1210));
  OR3_X1    g784(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n705), .B2(new_n706), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1210), .A2(new_n994), .A3(new_n1212), .ZN(G225));
  INV_X1    g787(.A(G225), .ZN(G308));
endmodule


