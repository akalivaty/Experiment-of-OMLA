//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT74), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT28), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n220), .B1(new_n223), .B2(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT71), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n219), .C1(new_n225), .C2(new_n228), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT28), .A3(new_n227), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT72), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n233), .A2(new_n236), .A3(KEYINPUT28), .A4(new_n227), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n230), .A2(new_n232), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n218), .B1(new_n238), .B2(KEYINPUT73), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n237), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n227), .B(new_n226), .C1(new_n233), .C2(new_n220), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n231), .B1(new_n241), .B2(new_n219), .ZN(new_n242));
  INV_X1    g041(.A(new_n232), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n248), .A2(new_n249), .B1(new_n213), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT66), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n254), .B(KEYINPUT64), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n252), .A4(new_n251), .ZN(new_n260));
  NOR2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(KEYINPUT23), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n210), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n264), .A2(new_n268), .A3(new_n265), .A4(new_n210), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n257), .A2(new_n260), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n210), .B(KEYINPUT68), .Z(new_n273));
  NAND3_X1  g072(.A1(new_n205), .A2(KEYINPUT23), .A3(new_n207), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n213), .A2(new_n250), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n254), .C1(G183gat), .C2(G190gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n271), .B1(new_n262), .B2(new_n263), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n273), .A2(new_n274), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT29), .B1(new_n247), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n281), .B(KEYINPUT82), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n278), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n270), .B2(new_n271), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(new_n239), .B2(new_n246), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n280), .A2(new_n282), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G211gat), .ZN(new_n289));
  INV_X1    g088(.A(G218gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n296), .A2(KEYINPUT81), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT81), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(KEYINPUT81), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n292), .A3(new_n291), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT92), .B1(new_n288), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n284), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT83), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n215), .A2(new_n217), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT73), .B(new_n240), .C1(new_n242), .C2(new_n243), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n238), .A2(KEYINPUT73), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n279), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n284), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n282), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n308), .A2(new_n304), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n287), .A2(new_n281), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n307), .B2(KEYINPUT83), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT92), .A3(new_n304), .A4(new_n317), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT37), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT93), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT38), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n319), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT93), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT37), .A4(new_n323), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  AOI221_X4 g131(.A(new_n305), .B1(new_n313), .B2(new_n283), .C1(new_n315), .C2(new_n281), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n308), .A2(new_n317), .A3(new_n318), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(new_n305), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT37), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n325), .A2(new_n326), .A3(new_n329), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n332), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n283), .B1(new_n313), .B2(new_n314), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n318), .B1(new_n340), .B2(new_n316), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n307), .A2(KEYINPUT83), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n305), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n333), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n339), .B1(new_n345), .B2(KEYINPUT37), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n335), .A2(new_n336), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT38), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n332), .A3(new_n344), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  INV_X1    g149(.A(G127gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(G134gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(G127gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT77), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G113gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .A4(G120gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT78), .B1(new_n356), .B2(G120gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT77), .B(G113gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(G120gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT79), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(new_n359), .A3(G120gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n363), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n361), .A4(new_n355), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT75), .A2(G134gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT75), .A2(G134gat), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(new_n351), .ZN(new_n375));
  OR3_X1    g174(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n354), .ZN(new_n376));
  XOR2_X1   g175(.A(G113gat), .B(G120gat), .Z(new_n377));
  AOI22_X1  g176(.A1(new_n375), .A2(KEYINPUT76), .B1(new_n377), .B2(new_n350), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT2), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(G155gat), .B2(G162gat), .ZN(new_n388));
  INV_X1    g187(.A(G141gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(G148gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT84), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n386), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n383), .B1(new_n387), .B2(new_n384), .ZN(new_n399));
  OR2_X1    g198(.A1(KEYINPUT85), .A2(G148gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT85), .A2(G148gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(G141gat), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n379), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n366), .A2(new_n371), .B1(new_n376), .B2(new_n378), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n398), .A2(KEYINPUT3), .A3(new_n403), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414));
  INV_X1    g213(.A(G155gat), .ZN(new_n415));
  INV_X1    g214(.A(G162gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT2), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n396), .B2(KEYINPUT84), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n393), .A2(new_n394), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n385), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n390), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n386), .A3(new_n417), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n412), .B1(new_n424), .B2(new_n380), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n410), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n404), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n380), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT86), .A3(new_n408), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n407), .A2(KEYINPUT86), .A3(new_n404), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n412), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(KEYINPUT5), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(new_n398), .B2(new_n403), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n420), .A2(new_n414), .A3(new_n422), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n411), .C1(new_n436), .C2(new_n407), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n407), .A2(KEYINPUT4), .A3(new_n404), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n379), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT80), .B1(new_n372), .B2(new_n379), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n440), .A2(new_n441), .A3(new_n427), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n438), .B(new_n439), .C1(new_n442), .C2(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n448), .A3(new_n443), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n451), .B(new_n448), .C1(new_n432), .C2(new_n443), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n349), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n338), .A2(new_n348), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n429), .A2(new_n430), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT39), .B1(new_n459), .B2(new_n412), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n424), .A2(new_n380), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(new_n439), .C1(new_n442), .C2(KEYINPUT4), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n412), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n464), .A3(new_n412), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n448), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(KEYINPUT90), .A3(new_n448), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT40), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n448), .B1(new_n432), .B2(new_n443), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n470), .B2(new_n473), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n335), .A2(new_n477), .A3(new_n332), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n304), .B1(new_n322), .B2(new_n317), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n339), .B1(new_n479), .B2(new_n333), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n349), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n474), .A2(new_n476), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n304), .B1(new_n314), .B2(new_n435), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT29), .B1(new_n301), .B2(new_n303), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n427), .B1(new_n486), .B2(KEYINPUT3), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n487), .B2(KEYINPUT87), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n427), .C1(new_n486), .C2(KEYINPUT3), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n427), .B(KEYINPUT88), .C1(new_n486), .C2(KEYINPUT3), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n305), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n484), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(G22gat), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  XNOR2_X1  g298(.A(G78gat), .B(G106gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT31), .B(G50gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n491), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n493), .A2(new_n496), .ZN(new_n504));
  INV_X1    g303(.A(G22gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n499), .A2(new_n502), .B1(new_n506), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n508), .A2(new_n506), .A3(new_n498), .A4(new_n502), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n458), .A2(new_n482), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n481), .A2(new_n478), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n453), .A2(new_n455), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n507), .A2(new_n509), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  XOR2_X1   g315(.A(G15gat), .B(G43gat), .Z(new_n517));
  XNOR2_X1  g316(.A(G71gat), .B(G99gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G227gat), .ZN(new_n521));
  INV_X1    g320(.A(G233gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n382), .A2(new_n405), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n313), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n440), .A2(new_n441), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n247), .B2(new_n279), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n313), .A2(new_n524), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n247), .A2(new_n526), .A3(new_n279), .ZN(new_n532));
  INV_X1    g331(.A(new_n523), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT34), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT34), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n531), .A2(new_n532), .A3(new_n536), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n532), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT33), .B1(new_n540), .B2(new_n523), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n535), .B(new_n537), .C1(new_n541), .C2(new_n520), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n528), .A2(KEYINPUT32), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n539), .B2(new_n542), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n516), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n543), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT36), .A3(new_n545), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n514), .A2(new_n515), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n511), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n510), .A2(new_n550), .A3(new_n545), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT35), .B1(new_n514), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n546), .A2(new_n515), .A3(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT35), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n452), .A2(new_n451), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n475), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n454), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n481), .B2(new_n478), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT41), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G29gat), .ZN(new_n570));
  INV_X1    g369(.A(G36gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT14), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT14), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n574), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G43gat), .B(G50gat), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n575), .A2(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n581), .A2(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n582), .B2(new_n587), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n585), .A2(KEYINPUT97), .A3(KEYINPUT17), .A4(new_n579), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT101), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n565), .A2(KEYINPUT41), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n586), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n603), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n606), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n569), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n607), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n568), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(KEYINPUT99), .ZN(new_n623));
  XOR2_X1   g422(.A(G57gat), .B(G64gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(KEYINPUT99), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G71gat), .B(G78gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G127gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G15gat), .B(G22gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(G1gat), .ZN(new_n636));
  OAI21_X1  g435(.A(G8gat), .B1(new_n636), .B2(KEYINPUT96), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT16), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(G1gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n638), .A2(new_n639), .A3(G1gat), .ZN(new_n642));
  OAI22_X1  g441(.A1(new_n641), .A2(new_n642), .B1(G1gat), .B2(new_n635), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n637), .B(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(new_n629), .B2(new_n630), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n634), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n415), .ZN(new_n648));
  XOR2_X1   g447(.A(G183gat), .B(G211gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n646), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n621), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G197gat), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT11), .B(G169gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n588), .A2(new_n644), .A3(new_n590), .A4(new_n591), .ZN(new_n659));
  NAND2_X1  g458(.A1(G229gat), .A2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n644), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n584), .A2(new_n586), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n658), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n660), .B(KEYINPUT13), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n610), .A2(new_n644), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n662), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n663), .B2(new_n664), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n659), .A2(KEYINPUT18), .A3(new_n660), .A4(new_n662), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT98), .B1(new_n663), .B2(new_n664), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(new_n673), .C1(new_n676), .C2(new_n658), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n603), .A2(new_n629), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n600), .A2(new_n602), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n600), .A2(new_n602), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n628), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n603), .A2(new_n629), .A3(KEYINPUT103), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT10), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n680), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n680), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n686), .A2(new_n692), .A3(new_n687), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(KEYINPUT105), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n691), .A2(new_n693), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT105), .B1(new_n694), .B2(new_n698), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n653), .A2(new_n679), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n564), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n560), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G1gat), .ZN(G1324gat));
  INV_X1    g507(.A(new_n512), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT16), .B(G8gat), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n706), .A2(new_n709), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n711), .A2(new_n712), .B1(new_n713), .B2(G8gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(new_n706), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n546), .A2(new_n547), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n720), .A2(G15gat), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n548), .A2(new_n551), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n515), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  AOI22_X1  g528(.A1(new_n511), .A2(new_n552), .B1(new_n555), .B2(new_n562), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n620), .ZN(new_n731));
  INV_X1    g530(.A(new_n651), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n679), .A3(new_n704), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n570), .A3(new_n560), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n730), .B2(new_n620), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n546), .A2(new_n547), .A3(new_n516), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT36), .B1(new_n550), .B2(new_n545), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n741), .A2(new_n742), .B1(new_n561), .B2(new_n510), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n345), .A2(KEYINPUT37), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n337), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n456), .B1(new_n745), .B2(KEYINPUT38), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n515), .B1(new_n746), .B2(new_n338), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n482), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n514), .A2(new_n554), .A3(KEYINPUT35), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n557), .B1(new_n556), .B2(new_n561), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT44), .B(new_n621), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n740), .A2(new_n752), .A3(new_n733), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n752), .A3(KEYINPUT109), .A4(new_n733), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n560), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n570), .B1(new_n757), .B2(KEYINPUT110), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT110), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n736), .A2(new_n737), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n738), .A2(new_n759), .A3(new_n760), .ZN(G1328gat));
  AOI21_X1  g560(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n734), .A2(new_n709), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n755), .A2(new_n709), .A3(new_n756), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n571), .B2(new_n766), .ZN(G1329gat));
  INV_X1    g566(.A(G43gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n734), .A2(new_n768), .A3(new_n721), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n724), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n772), .A3(new_n756), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(G43gat), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G43gat), .B1(new_n753), .B2(new_n724), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n770), .B1(new_n775), .B2(new_n769), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1330gat));
  OAI21_X1  g578(.A(G50gat), .B1(new_n753), .B2(new_n510), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n510), .A2(G50gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n734), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(KEYINPUT48), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n755), .A2(new_n515), .A3(new_n756), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G50gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n782), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n782), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n785), .B2(G50gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(KEYINPUT113), .A3(KEYINPUT48), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n783), .B1(new_n789), .B2(new_n792), .ZN(G1331gat));
  NAND2_X1  g592(.A1(new_n679), .A2(new_n704), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n730), .A2(new_n653), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n560), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g596(.A1(new_n795), .A2(new_n709), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n798), .B2(new_n799), .ZN(G1333gat));
  NAND2_X1  g601(.A1(new_n795), .A2(new_n772), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n722), .A2(G71gat), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(G71gat), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n795), .A2(new_n515), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT114), .B(G78gat), .Z(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1335gat));
  NAND2_X1  g608(.A1(new_n651), .A2(new_n679), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n730), .A2(new_n620), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(KEYINPUT115), .A3(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT115), .B1(new_n811), .B2(KEYINPUT51), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n597), .A3(new_n560), .A4(new_n704), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n740), .A2(new_n752), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n732), .A2(new_n794), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822), .B2(new_n513), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1336gat));
  NOR3_X1   g623(.A1(new_n512), .A2(new_n703), .A3(G92gat), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(new_n709), .A3(new_n821), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G92gat), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n813), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n811), .A2(KEYINPUT51), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n833), .A2(new_n825), .B1(G92gat), .B2(new_n827), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n826), .A2(new_n830), .B1(new_n834), .B2(new_n829), .ZN(G1337gat));
  NOR3_X1   g634(.A1(new_n722), .A2(G99gat), .A3(new_n703), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G99gat), .B1(new_n822), .B2(new_n724), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1338gat));
  NOR3_X1   g638(.A1(new_n510), .A2(new_n703), .A3(G106gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(new_n816), .B2(new_n817), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n515), .A3(new_n821), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n842), .B2(G106gat), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(G106gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n831), .B2(new_n832), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(new_n843), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n845), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(G1339gat));
  INV_X1    g653(.A(new_n691), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n697), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n688), .A2(new_n680), .A3(new_n690), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT54), .A3(new_n691), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT55), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n700), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(KEYINPUT55), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n857), .A2(new_n859), .A3(new_n865), .A4(KEYINPUT55), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n678), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n671), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n665), .A2(new_n658), .A3(new_n673), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n660), .B1(new_n659), .B2(new_n662), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n670), .A2(new_n662), .A3(new_n669), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n657), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n701), .B2(new_n702), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n621), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n615), .A2(new_n619), .A3(new_n873), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n651), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n652), .A2(new_n679), .A3(new_n703), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n513), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n709), .A2(new_n554), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT118), .Z(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n364), .A3(new_n678), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n515), .B1(new_n879), .B2(new_n880), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n709), .A2(new_n513), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n721), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G113gat), .B1(new_n888), .B2(new_n679), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1340gat));
  INV_X1    g689(.A(G120gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n891), .A3(new_n704), .ZN(new_n892));
  OAI21_X1  g691(.A(G120gat), .B1(new_n888), .B2(new_n703), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1341gat));
  OAI21_X1  g693(.A(G127gat), .B1(new_n888), .B2(new_n651), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n732), .A2(new_n351), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n883), .B2(new_n896), .ZN(G1342gat));
  OR4_X1    g696(.A1(new_n374), .A2(new_n883), .A3(new_n373), .A4(new_n620), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n888), .B2(new_n620), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G1343gat));
  NAND2_X1  g701(.A1(new_n879), .A2(new_n880), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n515), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n724), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n873), .B(new_n910), .C1(new_n701), .C2(new_n702), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n867), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n878), .B1(new_n912), .B2(new_n620), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(new_n732), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n510), .B1(new_n914), .B2(new_n880), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n907), .B(new_n678), .C1(new_n908), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G141gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n772), .A2(new_n510), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n881), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n709), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n679), .A2(G141gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n881), .A2(new_n512), .A3(new_n918), .A4(new_n923), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT120), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n916), .B2(G141gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n929), .B2(new_n925), .ZN(G1344gat));
  AOI21_X1  g729(.A(KEYINPUT59), .B1(new_n400), .B2(new_n401), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n907), .B1(new_n908), .B2(new_n915), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n703), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n651), .B1(new_n913), .B2(KEYINPUT122), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n936), .B(new_n878), .C1(new_n620), .C2(new_n912), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n880), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n510), .A2(KEYINPUT57), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n906), .A2(new_n703), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G148gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n934), .B1(new_n944), .B2(KEYINPUT59), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT123), .B(new_n946), .C1(new_n943), .C2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n933), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n922), .A2(new_n400), .A3(new_n401), .A4(new_n704), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1345gat));
  OAI21_X1  g749(.A(G155gat), .B1(new_n932), .B2(new_n651), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n922), .A2(new_n415), .A3(new_n732), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n932), .B2(new_n620), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n922), .A2(new_n416), .A3(new_n621), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n512), .A2(new_n560), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n958), .A2(new_n722), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n886), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(new_n203), .A3(new_n679), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n560), .B1(new_n879), .B2(new_n880), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n554), .A2(new_n512), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n678), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n961), .B1(new_n203), .B2(new_n966), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n965), .B2(new_n704), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n886), .A2(G176gat), .A3(new_n704), .A4(new_n959), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1349gat));
  OAI21_X1  g771(.A(G183gat), .B1(new_n960), .B2(new_n651), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n732), .A2(new_n233), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g775(.A(G190gat), .B1(new_n960), .B2(new_n620), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT61), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n965), .A2(new_n227), .A3(new_n621), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1351gat));
  NOR3_X1   g779(.A1(new_n772), .A2(new_n512), .A3(new_n510), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(G197gat), .B1(new_n983), .B2(new_n678), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n938), .A2(new_n939), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n772), .A2(new_n958), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n678), .A2(G197gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(G1352gat));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(G204gat), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n982), .A2(new_n703), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT62), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n991), .B1(new_n987), .B2(new_n703), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1353gat));
  NAND3_X1  g794(.A1(new_n983), .A2(new_n289), .A3(new_n732), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n940), .A2(new_n732), .A3(new_n941), .A4(new_n986), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n985), .A2(KEYINPUT126), .A3(new_n732), .A4(new_n986), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  AOI22_X1  g802(.A1(new_n1001), .A2(new_n1003), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n1004));
  NAND2_X1  g803(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1005));
  AOI211_X1 g804(.A(new_n1005), .B(new_n1002), .C1(new_n999), .C2(new_n1000), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n996), .B1(new_n1004), .B2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(G218gat), .B1(new_n987), .B2(new_n620), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n983), .A2(new_n290), .A3(new_n621), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1355gat));
endmodule


