//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n466), .B(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G137), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n483), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n482), .A2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND3_X1  g069(.A1(new_n463), .A2(G102), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n464), .B2(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(new_n463), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n479), .A2(new_n481), .A3(G138), .A4(new_n463), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .A4(new_n463), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT69), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n495), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n479), .A2(new_n481), .A3(G126), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n496), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n509), .A2(new_n510), .A3(new_n502), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n516), .A2(new_n518), .A3(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(G651), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(new_n525), .B1(new_n522), .B2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G50), .A3(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(G88), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n527), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n528), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(new_n525), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n522), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n534), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n533), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n538), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n524), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n516), .A2(new_n518), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n526), .A2(G81), .A3(new_n528), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT72), .B(G43), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n526), .A2(G543), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT73), .Z(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G188));
  NAND4_X1  g143(.A1(new_n535), .A2(G91), .A3(new_n536), .A4(new_n528), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n526), .A2(new_n571), .A3(G91), .A4(new_n528), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n517), .A2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT76), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G65), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n524), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n535), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n588), .ZN(G299));
  OAI21_X1  g164(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n526), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G49), .ZN(new_n592));
  INV_X1    g167(.A(G87), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n591), .B2(new_n592), .C1(new_n593), .C2(new_n532), .ZN(G288));
  NAND2_X1  g169(.A1(new_n533), .A2(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n538), .A2(G48), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n524), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n552), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n538), .A2(G47), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n533), .A2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT76), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT76), .B1(new_n516), .B2(new_n518), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT77), .B(G66), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT78), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n577), .A2(new_n578), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n611), .C1(new_n615), .C2(new_n609), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(G651), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n538), .A2(G54), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n526), .A2(G92), .A3(new_n528), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n606), .B1(new_n623), .B2(G868), .ZN(G284));
  XOR2_X1   g199(.A(G284), .B(KEYINPUT80), .Z(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  XOR2_X1   g201(.A(G299), .B(KEYINPUT81), .Z(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n476), .A2(new_n464), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR3_X1    g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n483), .A2(G135), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n645), .B(new_n646), .C1(G111), .C2(new_n463), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n489), .A2(G123), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n642), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  OAI21_X1  g225(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n639), .A2(new_n640), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n641), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n660), .A2(KEYINPUT16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n660), .A2(KEYINPUT16), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(KEYINPUT17), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n684), .B(new_n677), .C1(KEYINPUT17), .C2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(KEYINPUT87), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n678), .A2(KEYINPUT87), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT88), .Z(new_n690));
  XNOR2_X1  g265(.A(G2096), .B(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G227));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n703), .A2(new_n700), .A3(new_n698), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n698), .A2(new_n694), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n702), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n701), .B(new_n704), .C1(new_n706), .C2(new_n700), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT99), .B(G1966), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G11), .ZN(new_n719));
  INV_X1    g294(.A(G28), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n720), .B2(KEYINPUT30), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT30), .B2(new_n720), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT90), .A2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT90), .A2(G29), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n722), .B1(new_n649), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n729), .B2(G1961), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n718), .A2(new_n719), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G34), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n726), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n486), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n483), .A2(G139), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n463), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G2072), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n726), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n726), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT29), .B(G2090), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n748), .B(new_n752), .C1(G1961), .C2(new_n729), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n737), .A2(G32), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT97), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n476), .A2(G105), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n489), .A2(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n483), .A2(G141), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(new_n737), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT98), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n763), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n725), .A2(G27), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n725), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2078), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n741), .A2(new_n753), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G20), .ZN(new_n772));
  INV_X1    g347(.A(G299), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n714), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n772), .B(new_n774), .S(KEYINPUT23), .Z(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n770), .A2(new_n771), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n623), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n714), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n560), .B2(new_n714), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1341), .Z(new_n785));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n726), .B2(G26), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n726), .A2(KEYINPUT28), .A3(G26), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n483), .A2(G140), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  OR2_X1    g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n489), .A2(G128), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n786), .B(new_n788), .C1(new_n794), .C2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n782), .A2(new_n785), .A3(new_n796), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n732), .B(new_n778), .C1(KEYINPUT95), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n714), .A2(G24), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n603), .A2(new_n604), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n714), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1986), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n714), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n804));
  XNOR2_X1  g379(.A(G288), .B(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n803), .B1(new_n805), .B2(new_n714), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT33), .B(G1976), .Z(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n714), .A2(G6), .ZN(new_n809));
  INV_X1    g384(.A(G305), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n714), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n806), .A2(new_n807), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n714), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n714), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n808), .A2(new_n813), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n802), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n483), .A2(G131), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n489), .A2(G119), .ZN(new_n823));
  NOR2_X1   g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(new_n725), .Z(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G1991), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT91), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n821), .B(new_n830), .C1(new_n820), .C2(new_n819), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n738), .A2(new_n739), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n797), .A2(KEYINPUT95), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n798), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(G150));
  INV_X1    g411(.A(G150), .ZN(G311));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n552), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n538), .A2(G55), .B1(G651), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n533), .A2(G93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n623), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n555), .A2(new_n556), .A3(new_n558), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n841), .A2(new_n850), .A3(new_n842), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n559), .B2(KEYINPUT102), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n559), .A2(KEYINPUT102), .A3(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n851), .B1(new_n858), .B2(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n848), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n845), .B1(new_n862), .B2(G860), .ZN(G145));
  NAND2_X1  g438(.A1(new_n483), .A2(G142), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n489), .A2(G130), .ZN(new_n865));
  NOR2_X1   g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n746), .B(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n826), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n502), .A2(new_n503), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n502), .B2(new_n503), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n509), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n794), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n762), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n794), .A2(new_n877), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n876), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n762), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n882), .A2(new_n885), .A3(new_n637), .ZN(new_n886));
  INV_X1    g461(.A(new_n637), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n762), .A3(new_n878), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n871), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n637), .B1(new_n882), .B2(new_n885), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(new_n887), .A3(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n870), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n649), .B(new_n493), .Z(new_n897));
  XNOR2_X1  g472(.A(G160), .B(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n896), .ZN(new_n902));
  INV_X1    g477(.A(new_n898), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT105), .B(G37), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g483(.A(G288), .B(KEYINPUT93), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n800), .A2(G303), .ZN(new_n910));
  NAND2_X1  g485(.A1(G290), .A2(G166), .ZN(new_n911));
  AOI21_X1  g486(.A(G305), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(G305), .A3(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n916), .A2(new_n912), .A3(new_n805), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n632), .A2(new_n861), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n623), .A2(new_n630), .A3(new_n860), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n582), .B2(new_n588), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NOR4_X1   g502(.A1(new_n573), .A2(new_n587), .A3(new_n581), .A4(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n622), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n622), .A2(new_n927), .A3(G299), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT41), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n579), .A2(new_n580), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n570), .B(new_n572), .C1(new_n933), .C2(new_n524), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n934), .B2(new_n587), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n582), .A2(KEYINPUT107), .A3(new_n588), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n622), .A2(new_n927), .A3(G299), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n925), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n925), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n924), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n929), .A2(new_n930), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n922), .A2(new_n923), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n921), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n920), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT109), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n955), .A2(new_n943), .B1(new_n922), .B2(new_n923), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT108), .B1(new_n956), .B2(new_n949), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n918), .B(KEYINPUT42), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G868), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  INV_X1    g537(.A(G868), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n843), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n951), .B2(new_n959), .ZN(new_n966));
  INV_X1    g541(.A(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT110), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(G295));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n964), .ZN(G331));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n915), .B2(new_n917), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n805), .B1(new_n916), .B2(new_n912), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n913), .A2(new_n909), .A3(new_n914), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT112), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(G168), .A2(G301), .ZN(new_n977));
  NAND2_X1  g552(.A1(G171), .A2(G286), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n860), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n859), .A3(new_n857), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n955), .B2(new_n943), .ZN(new_n985));
  INV_X1    g560(.A(new_n946), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n987), .A3(new_n982), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n860), .A2(KEYINPUT111), .A3(new_n979), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n976), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n941), .B2(new_n944), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n946), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n994), .A3(new_n918), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  OR3_X1    g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n953), .A2(new_n954), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n993), .A2(new_n1000), .B1(new_n986), .B2(new_n983), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n905), .B1(new_n1001), .B2(new_n976), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n995), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n998), .B1(new_n997), .B2(KEYINPUT43), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n999), .A2(KEYINPUT44), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n997), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n997), .B2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1009), .A3(new_n995), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g588(.A1(new_n504), .A2(KEYINPUT104), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n873), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n1015), .B2(new_n509), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(KEYINPUT45), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n477), .A2(G40), .A3(new_n484), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n472), .A2(new_n1018), .A3(new_n473), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT115), .Z(new_n1021));
  INV_X1    g596(.A(G2067), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n883), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n794), .A2(G2067), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n762), .B(G1996), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n826), .A2(new_n828), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n826), .A2(new_n828), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1986), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n800), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G290), .A2(G1986), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1021), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n505), .A2(new_n511), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1019), .B(new_n1040), .C1(new_n1016), .C2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n876), .A2(new_n1039), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT50), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(KEYINPUT118), .A3(new_n1019), .A4(new_n1040), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n505), .A2(new_n511), .A3(new_n1039), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1039), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1019), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n817), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1037), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g634(.A(KEYINPUT116), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1049), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n876), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1044), .A3(new_n1065), .A4(new_n1019), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1037), .B(new_n1062), .C1(new_n1054), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n1055), .A2(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G2090), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1070), .A2(new_n1047), .B1(new_n817), .B2(new_n1053), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT119), .B(new_n1062), .C1(new_n1071), .C2(new_n1037), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT117), .B(G1981), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n810), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G305), .A2(G1981), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT49), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(G8), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n909), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n805), .A2(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(G8), .A3(new_n1079), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1064), .A2(new_n1019), .A3(new_n1065), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n505), .A2(new_n511), .A3(KEYINPUT45), .A4(new_n1039), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1019), .B(new_n1093), .C1(new_n1016), .C2(KEYINPUT45), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1092), .A2(new_n739), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n1037), .A3(G286), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1069), .A2(new_n1072), .A3(new_n1090), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1063), .B1(new_n1101), .B2(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1089), .B1(new_n1102), .B2(KEYINPUT119), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1103), .A2(KEYINPUT120), .A3(new_n1069), .A4(new_n1097), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1054), .A2(new_n1066), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1062), .B1(new_n1107), .B2(new_n1037), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(new_n1097), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1067), .A2(new_n1105), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1090), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1090), .A2(new_n1097), .A3(new_n1108), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1106), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1053), .B2(G2078), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1091), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1118), .A2(G2078), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1119), .B(new_n1121), .C1(new_n1094), .C2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(G301), .B(KEYINPUT54), .Z(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1069), .A2(new_n1072), .A3(new_n1090), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(G286), .A2(G8), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT51), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1128), .B(new_n1132), .C1(new_n1096), .C2(new_n1037), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G2084), .B2(new_n1091), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n1131), .C1(new_n1135), .C2(G286), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(G8), .A3(G286), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1121), .B(KEYINPUT126), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1052), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1017), .A2(new_n1140), .A3(new_n1122), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1018), .A2(new_n469), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1139), .A2(new_n1124), .A3(new_n1119), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1127), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1041), .A2(new_n776), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n582), .B2(KEYINPUT122), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G299), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n582), .B(new_n588), .C1(KEYINPUT122), .C2(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT123), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1051), .A2(new_n1019), .A3(new_n1052), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1147), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1091), .A2(new_n781), .ZN(new_n1156));
  INV_X1    g731(.A(new_n473), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(new_n471), .A3(G40), .A4(new_n485), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1045), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1022), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(new_n1161), .A3(new_n932), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1151), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1160), .A4(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1161), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1091), .A2(new_n781), .B1(new_n1159), .B2(new_n1022), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1167), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n1165), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1155), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1163), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1164), .A2(KEYINPUT61), .A3(new_n1155), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT58), .B(G1341), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1053), .A2(G1996), .B1(new_n1159), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT59), .B1(new_n1180), .B2(new_n560), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1162), .B(new_n1164), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1146), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(G288), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1081), .A2(new_n1082), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1084), .B1(new_n1187), .B2(new_n1074), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1067), .B2(new_n1090), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1069), .A2(new_n1072), .A3(new_n1090), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1123), .A2(G171), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1138), .A2(KEYINPUT62), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1133), .A2(new_n1136), .A3(new_n1193), .A4(new_n1137), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1189), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1036), .B1(new_n1117), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(G1996), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1021), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1025), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1021), .B1(new_n880), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1021), .A2(KEYINPUT46), .A3(new_n1198), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT47), .Z(new_n1206));
  NAND2_X1  g781(.A1(new_n1021), .A2(new_n1035), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n1207), .B(KEYINPUT48), .Z(new_n1208));
  AOI21_X1  g783(.A(new_n1208), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1023), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1021), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT127), .Z(new_n1212));
  NOR3_X1   g787(.A1(new_n1206), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1197), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1216));
  INV_X1    g790(.A(KEYINPUT113), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n997), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n1218), .A2(new_n1010), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G229), .A2(new_n461), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n672), .A2(new_n692), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n904), .B2(new_n906), .ZN(new_n1223));
  AND3_X1   g797(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(G308));
  NAND3_X1  g798(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(G225));
endmodule


