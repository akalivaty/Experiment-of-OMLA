//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n203), .A2(new_n204), .A3(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT92), .B(G8gat), .Z(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(G8gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT93), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n214), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G57gat), .B(G64gat), .Z(new_n218));
  INV_X1    g017(.A(G71gat), .ZN(new_n219));
  INV_X1    g018(.A(G78gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(KEYINPUT9), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G71gat), .B(G78gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n217), .B1(KEYINPUT21), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(KEYINPUT21), .ZN(new_n226));
  NAND2_X1  g025(.A1(G231gat), .A2(G233gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G127gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n225), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G155gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n230), .B(new_n234), .Z(new_n235));
  NAND2_X1  g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236));
  INV_X1    g035(.A(G85gat), .ZN(new_n237));
  INV_X1    g036(.A(G92gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(KEYINPUT8), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT99), .ZN(new_n240));
  NAND2_X1  g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT7), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G99gat), .B(G106gat), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(G29gat), .A2(G36gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT14), .ZN(new_n250));
  INV_X1    g049(.A(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT89), .B1(new_n251), .B2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G43gat), .B(G50gat), .Z(new_n258));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n250), .B(new_n257), .C1(KEYINPUT15), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(KEYINPUT15), .B2(new_n260), .ZN(new_n262));
  INV_X1    g061(.A(new_n258), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT15), .B(new_n263), .C1(new_n250), .C2(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT17), .B1(new_n265), .B2(KEYINPUT90), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n267), .B(new_n268), .C1(new_n262), .C2(new_n264), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n248), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n245), .A2(new_n247), .ZN(new_n271));
  AND2_X1   g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n265), .A2(new_n271), .B1(KEYINPUT41), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(KEYINPUT100), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n274), .B(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n279));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n278), .B(new_n281), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n235), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT102), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT101), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n247), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n224), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n248), .A2(new_n224), .A3(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI211_X1 g092(.A(KEYINPUT102), .B(KEYINPUT10), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(new_n298), .A3(new_n290), .ZN(new_n299));
  XNOR2_X1  g098(.A(G120gat), .B(G148gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G176gat), .B(G204gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT103), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n299), .ZN(new_n305));
  INV_X1    g104(.A(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n283), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(G197gat), .B(G204gat), .Z(new_n313));
  AOI21_X1  g112(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n311), .B(new_n316), .C1(KEYINPUT22), .C2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT27), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT27), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT28), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n337), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n344), .A2(KEYINPUT25), .A3(new_n346), .A4(new_n336), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT65), .ZN(new_n348));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT24), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(G183gat), .A3(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n348), .A3(new_n355), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n347), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(KEYINPUT64), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n344), .A2(new_n336), .A3(new_n346), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT25), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n343), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT70), .ZN(new_n369));
  AOI211_X1 g168(.A(KEYINPUT65), .B(new_n354), .C1(new_n350), .C2(new_n352), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT25), .B(new_n364), .C1(new_n356), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n364), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n343), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n369), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT26), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n335), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  AND2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n349), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT66), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n385));
  AOI221_X4 g184(.A(new_n379), .B1(new_n329), .B2(new_n330), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT67), .B1(new_n387), .B2(new_n331), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n375), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n369), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n378), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n369), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n343), .A2(new_n379), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(KEYINPUT67), .A3(new_n331), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n395), .A2(new_n396), .B1(new_n374), .B2(new_n371), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n321), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n367), .A2(new_n390), .A3(new_n377), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n394), .ZN(new_n402));
  INV_X1    g201(.A(new_n321), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n394), .C2(new_n397), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  AND3_X1   g206(.A1(new_n400), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n400), .B2(new_n404), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n408), .A2(KEYINPUT30), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n394), .B1(new_n412), .B2(new_n375), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n321), .B(new_n413), .C1(new_n401), .C2(new_n394), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n392), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n378), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n321), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT73), .B1(new_n418), .B2(new_n407), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n411), .B(new_n419), .C1(KEYINPUT30), .C2(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT83), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G106gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  XOR2_X1   g225(.A(G141gat), .B(G148gat), .Z(new_n427));
  INV_X1    g226(.A(G155gat), .ZN(new_n428));
  INV_X1    g227(.A(G162gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(KEYINPUT2), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G141gat), .B(G148gat), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n431), .B(new_n430), .C1(new_n435), .C2(KEYINPUT2), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n315), .A2(new_n438), .A3(new_n320), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n312), .B(KEYINPUT81), .C1(new_n313), .C2(new_n314), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n390), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n436), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n390), .B1(new_n444), .B2(KEYINPUT3), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n445), .A2(new_n321), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n426), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n321), .ZN(new_n448));
  INV_X1    g247(.A(new_n426), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n315), .B2(new_n320), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n444), .B1(new_n450), .B2(KEYINPUT3), .ZN(new_n451));
  AND4_X1   g250(.A1(KEYINPUT82), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n426), .B1(new_n445), .B2(new_n321), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT82), .B1(new_n453), .B2(new_n451), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n447), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G22gat), .ZN(new_n456));
  INV_X1    g255(.A(G22gat), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n447), .B(new_n457), .C1(new_n452), .C2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n220), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT80), .B(G78gat), .C1(new_n456), .C2(new_n458), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n425), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n458), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n453), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n457), .B1(new_n469), .B2(new_n447), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G78gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n459), .A2(new_n460), .A3(new_n220), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n424), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G120gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT1), .ZN(new_n477));
  XNOR2_X1  g276(.A(G127gat), .B(G134gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n389), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n478), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n477), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n412), .A2(new_n483), .A3(new_n375), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT34), .ZN(new_n486));
  XOR2_X1   g285(.A(G15gat), .B(G43gat), .Z(new_n487));
  XNOR2_X1  g286(.A(G71gat), .B(G99gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n480), .B2(new_n484), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(KEYINPUT33), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT32), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n480), .A2(new_n484), .ZN(new_n495));
  INV_X1    g294(.A(new_n481), .ZN(new_n496));
  AOI221_X4 g295(.A(new_n492), .B1(KEYINPUT33), .B2(new_n489), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n486), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  AOI221_X4 g297(.A(new_n479), .B1(new_n371), .B2(new_n374), .C1(new_n395), .C2(new_n396), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n483), .B1(new_n412), .B2(new_n375), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT32), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n489), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n485), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n489), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n501), .B(KEYINPUT32), .C1(new_n503), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n498), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n475), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n437), .A2(new_n442), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n444), .A2(KEYINPUT3), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n513), .A2(new_n514), .A3(new_n483), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g315(.A1(G225gat), .A2(G233gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT75), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT79), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n479), .B2(new_n444), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n479), .A2(new_n523), .A3(new_n444), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT79), .A3(new_n524), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n519), .A3(new_n524), .A4(new_n528), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n483), .B(new_n437), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n516), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G57gat), .B(G85gat), .Z(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G1gat), .B(G29gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(KEYINPUT6), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n536), .B2(KEYINPUT86), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(KEYINPUT86), .B2(new_n536), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n543), .A3(new_n535), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(KEYINPUT35), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n421), .A2(new_n512), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n507), .B1(new_n505), .B2(new_n509), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n559), .A3(new_n510), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(new_n475), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n400), .A2(new_n404), .ZN(new_n563));
  INV_X1    g362(.A(new_n407), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n410), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n404), .A4(new_n407), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n409), .A2(new_n410), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n565), .A4(new_n566), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n418), .A2(new_n407), .ZN(new_n572));
  INV_X1    g371(.A(new_n535), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n544), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n549), .A3(new_n550), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n571), .A2(new_n572), .B1(new_n576), .B2(new_n545), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n569), .A2(new_n570), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n555), .B(KEYINPUT35), .C1(new_n561), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n560), .A2(new_n475), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n570), .A2(new_n577), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n569), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n555), .B1(new_n583), .B2(KEYINPUT35), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n554), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n556), .A3(new_n559), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT69), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n511), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT69), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n586), .A2(new_n556), .A3(new_n559), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n570), .A2(new_n577), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT74), .B1(new_n411), .B2(new_n419), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n475), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT84), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n530), .A2(new_n515), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(KEYINPUT85), .A3(new_n518), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n513), .A2(new_n514), .A3(new_n483), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n527), .B2(new_n529), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n605), .B2(new_n519), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n533), .A2(new_n518), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n602), .A2(new_n606), .A3(KEYINPUT39), .A4(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n609), .A2(KEYINPUT40), .A3(new_n611), .A4(new_n543), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(new_n548), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n609), .A2(new_n543), .A3(new_n611), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n420), .B(new_n613), .C1(KEYINPUT40), .C2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n463), .A2(new_n474), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n407), .B1(new_n418), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n417), .A2(new_n403), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n402), .B1(new_n394), .B2(new_n397), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n619), .B(KEYINPUT37), .C1(new_n403), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT38), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n563), .B2(KEYINPUT37), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n552), .A2(new_n572), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n615), .B(new_n616), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n600), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n585), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G197gat), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT11), .B(G169gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  INV_X1    g433(.A(new_n265), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n216), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n213), .A2(new_n265), .A3(new_n215), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n217), .A2(new_n641), .A3(new_n265), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n216), .B1(new_n266), .B2(new_n269), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT94), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n216), .B(new_n647), .C1(new_n266), .C2(new_n269), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n646), .A2(new_n639), .A3(new_n637), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n648), .A2(new_n637), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n652), .A2(KEYINPUT18), .A3(new_n639), .A4(new_n646), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n634), .B1(new_n644), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n643), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n634), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n651), .A4(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(KEYINPUT97), .B(new_n634), .C1(new_n644), .C2(new_n654), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n310), .B1(new_n629), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT98), .B(new_n663), .C1(new_n585), .C2(new_n628), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n309), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n669), .B(new_n309), .C1(new_n665), .C2(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n576), .A2(new_n545), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(G8gat), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n671), .B2(new_n420), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n421), .B(new_n678), .C1(new_n668), .C2(new_n670), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT42), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n420), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n511), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n593), .B1(new_n668), .B2(new_n670), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n475), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n597), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n627), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n585), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n554), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT35), .B1(new_n561), .B2(new_n578), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT87), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(new_n579), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT106), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n585), .A2(new_n695), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n694), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n282), .A2(KEYINPUT44), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n282), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n629), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n308), .A2(new_n235), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n664), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n672), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n709), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n672), .A2(G29gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n719), .B(new_n720), .C1(new_n665), .C2(new_n666), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n717), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n714), .B1(new_n708), .B2(new_n711), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n251), .B1(new_n727), .B2(new_n673), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT107), .B1(new_n728), .B2(new_n723), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1328gat));
  OAI21_X1  g529(.A(G36gat), .B1(new_n716), .B2(new_n421), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n421), .A2(G36gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n719), .B(new_n732), .C1(new_n665), .C2(new_n666), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n252), .B1(new_n727), .B2(new_n420), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT108), .B1(new_n738), .B2(new_n734), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n593), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n712), .A2(G43gat), .A3(new_n741), .A4(new_n715), .ZN(new_n742));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n629), .A2(new_n664), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n629), .A2(new_n310), .A3(new_n664), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n719), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n748), .B2(new_n511), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n742), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n742), .A2(new_n750), .A3(new_n749), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n751), .ZN(G1330gat));
  NAND2_X1  g553(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n718), .B1(new_n745), .B2(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n616), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(G50gat), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G50gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n616), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n727), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT48), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n757), .A3(new_n719), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n475), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n756), .A2(new_n757), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n727), .A2(new_n761), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(new_n770), .ZN(G1331gat));
  AND2_X1   g570(.A1(new_n702), .A2(new_n706), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n664), .A2(new_n283), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n308), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n672), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n421), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT49), .B(G64gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n779), .B2(new_n782), .ZN(G1333gat));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n741), .A3(new_n775), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G71gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n686), .A2(new_n219), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n776), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n785), .B(KEYINPUT50), .C1(new_n776), .C2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1334gat));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n616), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT112), .B(G78gat), .Z(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1335gat));
  INV_X1    g593(.A(new_n235), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n663), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n308), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n708), .B2(new_n711), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n672), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n696), .A2(new_n701), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n796), .A2(new_n282), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT51), .B(new_n804), .C1(new_n696), .C2(new_n701), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(KEYINPUT113), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n802), .C1(new_n803), .C2(new_n805), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n308), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n673), .A2(new_n237), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n801), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  AOI21_X1  g612(.A(new_n238), .B1(new_n799), .B2(new_n420), .ZN(new_n814));
  INV_X1    g613(.A(new_n308), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(G92gat), .A3(new_n421), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n806), .B2(new_n807), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n808), .A2(new_n810), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n817), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n814), .B2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n800), .B2(new_n593), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n511), .A2(G99gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n811), .B2(new_n825), .ZN(G1338gat));
  INV_X1    g625(.A(G106gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n799), .B2(new_n475), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n308), .A2(new_n827), .A3(new_n475), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT114), .Z(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n806), .B2(new_n807), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT53), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n821), .B2(new_n830), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n828), .B2(new_n834), .ZN(G1339gat));
  NAND2_X1  g634(.A1(new_n773), .A2(new_n815), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n652), .A2(new_n646), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n640), .B1(new_n638), .B2(new_n642), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n837), .A2(new_n639), .B1(KEYINPUT115), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n633), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n659), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n297), .A2(KEYINPUT54), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n298), .B(new_n284), .C1(new_n293), .C2(new_n294), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n297), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n306), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n306), .A4(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n304), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n842), .A2(new_n850), .A3(new_n282), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n308), .A2(new_n841), .A3(new_n659), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n663), .B2(new_n850), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(new_n282), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n836), .B1(new_n854), .B2(new_n235), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n421), .A2(new_n673), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(new_n581), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(G113gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n664), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n512), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n856), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n512), .A4(new_n857), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n664), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(new_n866), .A3(G113gat), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n865), .B2(G113gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  AOI21_X1  g668(.A(G120gat), .B1(new_n858), .B2(new_n308), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n863), .A2(new_n864), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n308), .A2(G120gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1341gat));
  NAND3_X1  g672(.A1(new_n863), .A2(new_n235), .A3(new_n864), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G127gat), .ZN(new_n875));
  INV_X1    g674(.A(G127gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n876), .A3(new_n235), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1342gat));
  NOR2_X1   g681(.A1(new_n282), .A2(G134gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT121), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n887), .A3(KEYINPUT56), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n884), .B2(KEYINPUT56), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n891), .A4(new_n883), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n886), .A2(new_n888), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n863), .A2(new_n709), .A3(new_n864), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT120), .B1(new_n894), .B2(G134gat), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n894), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n741), .A2(new_n856), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT122), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n616), .A2(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n855), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n850), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n848), .A2(new_n304), .A3(KEYINPUT123), .A4(new_n849), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n903), .A2(new_n662), .A3(new_n661), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n709), .B1(new_n905), .B2(new_n852), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n795), .B1(new_n906), .B2(new_n851), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n616), .B1(new_n907), .B2(new_n836), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n901), .B(new_n664), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT124), .B1(new_n910), .B2(G141gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n741), .A2(new_n616), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n663), .A2(G141gat), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n857), .A2(new_n855), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n910), .B2(G141gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT58), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  AOI221_X4 g716(.A(new_n914), .B1(KEYINPUT124), .B2(new_n917), .C1(new_n910), .C2(G141gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(G1344gat));
  NOR2_X1   g718(.A1(new_n908), .A2(KEYINPUT57), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n855), .A2(KEYINPUT57), .A3(new_n475), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n899), .A2(new_n815), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n855), .A2(new_n857), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n912), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n308), .A2(new_n926), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n929), .A2(KEYINPUT125), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT125), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n924), .A2(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n934));
  OAI21_X1  g733(.A(G148gat), .B1(new_n934), .B2(new_n815), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n925), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1345gat));
  OAI21_X1  g736(.A(G155gat), .B1(new_n934), .B2(new_n795), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n235), .A2(new_n428), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n929), .B2(new_n939), .ZN(G1346gat));
  NOR3_X1   g739(.A1(new_n934), .A2(new_n429), .A3(new_n282), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n928), .A2(new_n709), .A3(new_n912), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n429), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n421), .A2(new_n673), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n855), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(new_n581), .ZN(new_n946));
  AOI21_X1  g745(.A(G169gat), .B1(new_n946), .B2(new_n664), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n944), .B(KEYINPUT126), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n862), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n332), .A3(new_n663), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n947), .A2(new_n950), .ZN(G1348gat));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n333), .A3(new_n308), .ZN(new_n952));
  OAI21_X1  g751(.A(G176gat), .B1(new_n949), .B2(new_n815), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  AND2_X1   g753(.A1(new_n323), .A2(new_n325), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n946), .A2(new_n955), .A3(new_n235), .ZN(new_n956));
  OAI21_X1  g755(.A(G183gat), .B1(new_n949), .B2(new_n795), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n949), .B2(new_n282), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT61), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n326), .A3(new_n709), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n741), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n922), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(G197gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n663), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n945), .A2(new_n912), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n945), .A2(new_n971), .A3(new_n912), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n664), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n966), .A2(new_n968), .B1(new_n973), .B2(new_n967), .ZN(G1352gat));
  OAI21_X1  g773(.A(G204gat), .B1(new_n965), .B2(new_n815), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n969), .A2(G204gat), .A3(new_n815), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  AND2_X1   g777(.A1(new_n970), .A2(new_n972), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n317), .A3(new_n235), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n235), .B(new_n964), .C1(new_n920), .C2(new_n921), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n965), .B2(new_n282), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n979), .A2(new_n318), .A3(new_n709), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


