

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U319 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n355) );
  XNOR2_X1 U320 ( .A(n356), .B(n355), .ZN(n393) );
  XNOR2_X1 U321 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U322 ( .A(n404), .B(KEYINPUT64), .ZN(n405) );
  XNOR2_X1 U323 ( .A(n327), .B(n326), .ZN(n331) );
  XNOR2_X1 U324 ( .A(n406), .B(n405), .ZN(n522) );
  NOR2_X1 U325 ( .A1(n430), .A2(n511), .ZN(n567) );
  XNOR2_X1 U326 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n288) );
  XNOR2_X1 U329 ( .A(G197GAT), .B(G211GAT), .ZN(n287) );
  XNOR2_X1 U330 ( .A(n288), .B(n287), .ZN(n306) );
  XNOR2_X1 U331 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n289), .B(KEYINPUT2), .ZN(n421) );
  XNOR2_X1 U333 ( .A(n306), .B(n421), .ZN(n303) );
  XOR2_X1 U334 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n291) );
  XNOR2_X1 U335 ( .A(KEYINPUT85), .B(KEYINPUT22), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U337 ( .A(G106GAT), .B(G148GAT), .Z(n359) );
  XOR2_X1 U338 ( .A(n359), .B(G204GAT), .Z(n293) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n342) );
  XNOR2_X1 U340 ( .A(n342), .B(G218GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U342 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U343 ( .A1(G228GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n298), .B(KEYINPUT86), .Z(n301) );
  XNOR2_X1 U346 ( .A(G22GAT), .B(G78GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n299), .B(G155GAT), .ZN(n333) );
  XNOR2_X1 U348 ( .A(n333), .B(KEYINPUT24), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n461) );
  XOR2_X1 U351 ( .A(G64GAT), .B(G204GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(G176GAT), .B(G92GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n364) );
  XNOR2_X1 U354 ( .A(n364), .B(n306), .ZN(n316) );
  XOR2_X1 U355 ( .A(G8GAT), .B(G183GAT), .Z(n320) );
  XOR2_X1 U356 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n311) );
  XOR2_X1 U357 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n308) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n440) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n309), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U362 ( .A(n440), .B(n341), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U364 ( .A(n320), .B(n312), .Z(n314) );
  NAND2_X1 U365 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n513) );
  INV_X1 U368 ( .A(KEYINPUT113), .ZN(n395) );
  XOR2_X1 U369 ( .A(G211GAT), .B(KEYINPUT77), .Z(n318) );
  XNOR2_X1 U370 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n322) );
  NAND2_X1 U373 ( .A1(G231GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(G57GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n323), .B(KEYINPUT13), .ZN(n363) );
  XNOR2_X1 U377 ( .A(n363), .B(KEYINPUT12), .ZN(n325) );
  INV_X1 U378 ( .A(KEYINPUT15), .ZN(n324) );
  XOR2_X1 U379 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n329) );
  XNOR2_X1 U380 ( .A(G127GAT), .B(KEYINPUT14), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(G15GAT), .ZN(n380) );
  XNOR2_X1 U385 ( .A(n380), .B(n333), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n548) );
  XOR2_X1 U387 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n337) );
  XNOR2_X1 U388 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n338), .B(G92GAT), .ZN(n340) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XOR2_X1 U392 ( .A(n367), .B(G106GAT), .Z(n339) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U394 ( .A(n342), .B(n341), .Z(n344) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n354) );
  XOR2_X1 U398 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n348) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G29GAT), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U401 ( .A(KEYINPUT70), .B(n349), .Z(n387) );
  XOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n351) );
  XNOR2_X1 U403 ( .A(G134GAT), .B(KEYINPUT67), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n387), .B(n352), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n538) );
  XOR2_X1 U407 ( .A(n538), .B(KEYINPUT36), .Z(n580) );
  NAND2_X1 U408 ( .A1(n548), .A2(n580), .ZN(n356) );
  XOR2_X1 U409 ( .A(G78GAT), .B(KEYINPUT32), .Z(n358) );
  XNOR2_X1 U410 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n357) );
  XOR2_X1 U411 ( .A(n358), .B(n357), .Z(n362) );
  XNOR2_X1 U412 ( .A(n359), .B(KEYINPUT33), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n360), .B(KEYINPUT31), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n366) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U417 ( .A(n368), .B(n367), .ZN(n370) );
  AND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U419 ( .A(n370), .B(n369), .ZN(n396) );
  XOR2_X1 U420 ( .A(G197GAT), .B(KEYINPUT69), .Z(n372) );
  XNOR2_X1 U421 ( .A(KEYINPUT68), .B(G141GAT), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n391) );
  XOR2_X1 U423 ( .A(G8GAT), .B(KEYINPUT29), .Z(n374) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(G36GAT), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U426 ( .A(G113GAT), .B(KEYINPUT72), .Z(n376) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(KEYINPUT30), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U429 ( .A(n378), .B(n377), .Z(n389) );
  INV_X1 U430 ( .A(n380), .ZN(n379) );
  NAND2_X1 U431 ( .A1(G169GAT), .A2(n379), .ZN(n383) );
  INV_X1 U432 ( .A(G169GAT), .ZN(n381) );
  NAND2_X1 U433 ( .A1(n381), .A2(n380), .ZN(n382) );
  NAND2_X1 U434 ( .A1(n383), .A2(n382), .ZN(n385) );
  NAND2_X1 U435 ( .A1(G229GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U437 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U438 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U439 ( .A(n391), .B(n390), .Z(n568) );
  NAND2_X1 U440 ( .A1(n396), .A2(n568), .ZN(n392) );
  NOR2_X1 U441 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U442 ( .A(n395), .B(n394), .ZN(n403) );
  XNOR2_X1 U443 ( .A(KEYINPUT111), .B(n548), .ZN(n563) );
  NAND2_X1 U444 ( .A1(n538), .A2(n563), .ZN(n400) );
  XNOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n398) );
  XNOR2_X1 U446 ( .A(KEYINPUT41), .B(n396), .ZN(n557) );
  INV_X1 U447 ( .A(n568), .ZN(n554) );
  NAND2_X1 U448 ( .A1(n557), .A2(n554), .ZN(n397) );
  XOR2_X1 U449 ( .A(n398), .B(n397), .Z(n399) );
  NOR2_X1 U450 ( .A1(n400), .A2(n399), .ZN(n401) );
  XOR2_X1 U451 ( .A(n401), .B(KEYINPUT47), .Z(n402) );
  NOR2_X1 U452 ( .A1(n403), .A2(n402), .ZN(n406) );
  XOR2_X1 U453 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n404) );
  NAND2_X1 U454 ( .A1(n513), .A2(n522), .ZN(n407) );
  XNOR2_X1 U455 ( .A(n407), .B(KEYINPUT54), .ZN(n430) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U457 ( .A(G1GAT), .B(G85GAT), .ZN(n408) );
  XNOR2_X1 U458 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U459 ( .A(G29GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U460 ( .A(n411), .B(n410), .ZN(n427) );
  XOR2_X1 U461 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n413) );
  XNOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n412) );
  XNOR2_X1 U463 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n415) );
  XNOR2_X1 U465 ( .A(G155GAT), .B(KEYINPUT1), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U467 ( .A(n417), .B(n416), .ZN(n425) );
  XOR2_X1 U468 ( .A(KEYINPUT89), .B(KEYINPUT93), .Z(n423) );
  XOR2_X1 U469 ( .A(G120GAT), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U470 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U472 ( .A(G113GAT), .B(n420), .Z(n444) );
  XNOR2_X1 U473 ( .A(n444), .B(n421), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n429) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n429), .B(n428), .ZN(n511) );
  NAND2_X1 U479 ( .A1(n461), .A2(n567), .ZN(n431) );
  XNOR2_X1 U480 ( .A(n431), .B(KEYINPUT55), .ZN(n449) );
  XOR2_X1 U481 ( .A(KEYINPUT65), .B(KEYINPUT83), .Z(n433) );
  XNOR2_X1 U482 ( .A(KEYINPUT81), .B(KEYINPUT84), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n448) );
  XOR2_X1 U484 ( .A(G176GAT), .B(G99GAT), .Z(n435) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U487 ( .A(KEYINPUT20), .B(G183GAT), .Z(n437) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(G71GAT), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U490 ( .A(n439), .B(n438), .Z(n446) );
  XOR2_X1 U491 ( .A(n440), .B(KEYINPUT82), .Z(n442) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U496 ( .A(n448), .B(n447), .ZN(n526) );
  NAND2_X1 U497 ( .A1(n449), .A2(n526), .ZN(n450) );
  XNOR2_X1 U498 ( .A(n450), .B(KEYINPUT121), .ZN(n558) );
  INV_X1 U499 ( .A(n558), .ZN(n562) );
  NOR2_X1 U500 ( .A1(n562), .A2(n538), .ZN(n454) );
  XNOR2_X1 U501 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n452) );
  INV_X1 U502 ( .A(G190GAT), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n472) );
  NAND2_X1 U504 ( .A1(n396), .A2(n554), .ZN(n486) );
  INV_X1 U505 ( .A(n538), .ZN(n551) );
  INV_X1 U506 ( .A(n548), .ZN(n577) );
  NOR2_X1 U507 ( .A1(n551), .A2(n577), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n455), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U509 ( .A(n461), .B(KEYINPUT28), .ZN(n525) );
  INV_X1 U510 ( .A(n525), .ZN(n517) );
  NOR2_X1 U511 ( .A1(n517), .A2(n526), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n513), .B(KEYINPUT27), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n459), .A2(n511), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT96), .B(n456), .Z(n523) );
  NAND2_X1 U515 ( .A1(n457), .A2(n523), .ZN(n468) );
  NOR2_X1 U516 ( .A1(n461), .A2(n526), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT26), .B(n458), .Z(n542) );
  INV_X1 U518 ( .A(n542), .ZN(n566) );
  NAND2_X1 U519 ( .A1(n566), .A2(n459), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n513), .A2(n526), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n462), .Z(n463) );
  NAND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n466) );
  INV_X1 U524 ( .A(n511), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n482) );
  NAND2_X1 U527 ( .A1(n469), .A2(n482), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT97), .B(n470), .Z(n501) );
  NOR2_X1 U529 ( .A1(n486), .A2(n501), .ZN(n479) );
  NAND2_X1 U530 ( .A1(n479), .A2(n511), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U532 ( .A(G1GAT), .B(n473), .Z(G1324GAT) );
  NAND2_X1 U533 ( .A1(n479), .A2(n513), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n476) );
  NAND2_X1 U536 ( .A1(n479), .A2(n526), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n478) );
  XOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT99), .Z(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XOR2_X1 U540 ( .A(G22GAT), .B(KEYINPUT101), .Z(n481) );
  NAND2_X1 U541 ( .A1(n479), .A2(n517), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n580), .A2(n482), .ZN(n483) );
  NOR2_X1 U544 ( .A1(n548), .A2(n483), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT103), .B(n484), .Z(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n485), .ZN(n510) );
  NOR2_X1 U547 ( .A1(n486), .A2(n510), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT38), .ZN(n498) );
  NAND2_X1 U549 ( .A1(n498), .A2(n511), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT105), .Z(n493) );
  NAND2_X1 U555 ( .A1(n513), .A2(n498), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n497) );
  XOR2_X1 U558 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n495) );
  NAND2_X1 U559 ( .A1(n498), .A2(n526), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n517), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  NAND2_X1 U566 ( .A1(n568), .A2(n557), .ZN(n509) );
  NOR2_X1 U567 ( .A1(n501), .A2(n509), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n511), .A2(n506), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n506), .A2(n513), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n526), .A2(n506), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U575 ( .A1(n506), .A2(n517), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n511), .A2(n518), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U583 ( .A1(n518), .A2(n526), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U588 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n529) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT115), .B(n524), .Z(n541) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n541), .A2(n527), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n533), .A2(n554), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U598 ( .A1(n533), .A2(n557), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  INV_X1 U600 ( .A(n533), .ZN(n537) );
  NOR2_X1 U601 ( .A1(n563), .A2(n537), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n554), .A2(n552), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U612 ( .A1(n552), .A2(n557), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT119), .Z(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n552), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U632 ( .A1(n568), .A2(n579), .ZN(n573) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT59), .B(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n396), .A2(n579), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  INV_X1 U644 ( .A(n579), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

