//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n206), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT72), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219));
  INV_X1    g018(.A(G211gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n215), .A2(new_n222), .A3(new_n218), .A4(new_n216), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n209), .ZN(new_n231));
  XNOR2_X1  g030(.A(G141gat), .B(G148gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(KEYINPUT2), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n224), .A2(new_n226), .B1(new_n225), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238));
  OR3_X1    g037(.A1(new_n229), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n213), .B1(new_n227), .B2(new_n235), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n240), .B2(new_n237), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT87), .B(G22gat), .Z(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT31), .B(G50gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n241), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(G22gat), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n246), .B(KEYINPUT86), .Z(new_n250));
  INV_X1    g049(.A(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(new_n243), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(G120gat), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(new_n258), .B2(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n256), .A3(G120gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G134gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G127gat), .ZN(new_n265));
  INV_X1    g064(.A(G127gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n256), .A2(G120gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n258), .A2(G113gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n270), .A2(new_n275), .A3(new_n233), .A4(new_n234), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n263), .A2(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n213), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT83), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n270), .A2(new_n275), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n278), .A2(KEYINPUT78), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT3), .B1(new_n211), .B2(new_n212), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n236), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n282), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT80), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT39), .ZN(new_n295));
  XOR2_X1   g094(.A(G1gat), .B(G29gat), .Z(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G57gat), .B(G85gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n213), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n276), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT39), .B1(new_n305), .B2(new_n293), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n294), .B1(new_n306), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT40), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n302), .B(KEYINPUT40), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT5), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n305), .B2(new_n293), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n293), .B1(new_n277), .B2(new_n280), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n317), .A2(KEYINPUT81), .A3(new_n290), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT81), .B1(new_n317), .B2(new_n290), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n282), .A2(new_n284), .A3(new_n290), .A4(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n301), .B1(new_n323), .B2(KEYINPUT89), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n320), .A2(KEYINPUT89), .A3(new_n322), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n224), .A2(new_n226), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT27), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT67), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT67), .B1(new_n333), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT28), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  INV_X1    g140(.A(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT26), .ZN(new_n343));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT26), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n343), .B(new_n344), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT66), .B1(new_n334), .B2(KEYINPUT27), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n332), .A3(G183gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT27), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n349), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT23), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n359), .A2(new_n361), .A3(new_n347), .ZN(new_n362));
  NAND3_X1  g161(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n334), .A2(new_n331), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n368), .A2(new_n363), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n331), .A3(new_n356), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT25), .A3(new_n362), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n340), .A2(new_n358), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT73), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n330), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n334), .A2(KEYINPUT27), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n332), .A2(G183gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n336), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n388), .B2(new_n331), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n346), .A2(new_n348), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n343), .A2(new_n344), .ZN(new_n391));
  INV_X1    g190(.A(new_n357), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT25), .B1(new_n362), .B2(new_n370), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT25), .A4(new_n347), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n375), .B2(new_n374), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n389), .A2(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n382), .B1(new_n398), .B2(new_n225), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n328), .B1(new_n381), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n380), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n329), .B1(new_n398), .B2(new_n382), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT75), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n373), .A2(new_n377), .ZN(new_n406));
  AOI21_X1  g205(.A(G190gat), .B1(new_n387), .B2(new_n336), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n358), .B1(new_n407), .B2(new_n383), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n380), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n405), .A2(new_n409), .B1(new_n410), .B2(new_n382), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n378), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n329), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n404), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n413), .A3(new_n420), .A4(new_n416), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n381), .A2(new_n399), .A3(new_n328), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT75), .B1(new_n401), .B2(new_n402), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n405), .B1(new_n398), .B2(new_n382), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n399), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n412), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n330), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n413), .A3(KEYINPUT76), .ZN(new_n432));
  INV_X1    g231(.A(new_n416), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n417), .A2(new_n419), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n422), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n254), .B1(new_n327), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n426), .A2(new_n430), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n431), .A2(KEYINPUT37), .A3(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n433), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(KEYINPUT91), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT91), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n446), .A3(new_n433), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n330), .B1(new_n411), .B2(new_n412), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n329), .B1(new_n378), .B2(new_n380), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(KEYINPUT37), .C1(new_n399), .C2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n439), .A3(new_n433), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n454), .B(new_n300), .C1(new_n320), .C2(new_n322), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n322), .A2(new_n300), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT6), .B1(new_n320), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n324), .B2(new_n325), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n418), .A2(new_n421), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n456), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n438), .B1(new_n448), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT71), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n378), .A2(new_n285), .ZN(new_n464));
  INV_X1    g263(.A(G227gat), .ZN(new_n465));
  INV_X1    g264(.A(G233gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n398), .A2(new_n278), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT32), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G15gat), .B(G43gat), .Z(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n475), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n469), .B(KEYINPUT32), .C1(new_n471), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n468), .ZN(new_n480));
  INV_X1    g279(.A(new_n467), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT34), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n485), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n476), .A3(new_n478), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n463), .B1(new_n490), .B2(KEYINPUT36), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n488), .A2(new_n493), .B1(new_n476), .B2(new_n478), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT36), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n487), .A2(KEYINPUT71), .A3(new_n496), .A4(new_n489), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n320), .A2(new_n322), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n458), .A2(new_n500), .B1(new_n501), .B2(new_n301), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n322), .A2(new_n300), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  INV_X1    g303(.A(new_n293), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n279), .B1(new_n213), .B2(new_n278), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n283), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n289), .A2(new_n236), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT78), .B1(new_n270), .B2(new_n275), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n270), .A2(KEYINPUT78), .A3(new_n275), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n504), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n317), .A2(KEYINPUT81), .A3(new_n290), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n514), .B2(new_n316), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT84), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n455), .B1(new_n502), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n499), .B1(new_n437), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n320), .A2(new_n457), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n500), .A3(new_n454), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n301), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n456), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n404), .A2(new_n413), .A3(KEYINPUT76), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT76), .B1(new_n404), .B2(new_n413), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n435), .B1(new_n526), .B2(new_n433), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(new_n527), .A3(KEYINPUT85), .A4(new_n422), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n498), .B1(new_n529), .B2(new_n254), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n492), .A2(new_n494), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n254), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n518), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n534));
  INV_X1    g333(.A(new_n490), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n254), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n459), .A2(new_n456), .ZN(new_n537));
  INV_X1    g336(.A(new_n437), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n462), .A2(new_n530), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n547));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT95), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT93), .B(G29gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n543), .B2(KEYINPUT15), .ZN(new_n556));
  INV_X1    g355(.A(G29gat), .ZN(new_n557));
  INV_X1    g356(.A(G36gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT14), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(G29gat), .B2(G36gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n554), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n551), .A2(new_n564), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n562), .A2(KEYINPUT92), .B1(new_n552), .B2(new_n558), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(KEYINPUT92), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n544), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n542), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n571), .A2(G1gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  INV_X1    g373(.A(G8gat), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(KEYINPUT96), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(KEYINPUT96), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n572), .A2(new_n574), .A3(new_n579), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n568), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT15), .B(new_n543), .C1(new_n582), .C2(new_n566), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n583), .B(KEYINPUT17), .C1(new_n564), .C2(new_n551), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n570), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n583), .B1(new_n564), .B2(new_n551), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n578), .A3(new_n580), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT18), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT18), .A4(new_n586), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n581), .B(new_n583), .C1(new_n564), .C2(new_n551), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n586), .B(KEYINPUT13), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G197gat), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT11), .B(G169gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n591), .A2(new_n602), .A3(new_n592), .A4(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n541), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G57gat), .B(G64gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT97), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G71gat), .B(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n610), .ZN(new_n615));
  OR2_X1    g414(.A1(G57gat), .A2(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(G57gat), .A2(G64gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT97), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT20), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n581), .B1(new_n622), .B2(new_n621), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G183gat), .B(G211gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n628), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G99gat), .A2(G106gat), .ZN(new_n636));
  INV_X1    g435(.A(G85gat), .ZN(new_n637));
  INV_X1    g436(.A(G92gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(KEYINPUT8), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT7), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G99gat), .B(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n642), .A2(new_n643), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n587), .A2(new_n650), .B1(KEYINPUT41), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n570), .B1(new_n647), .B2(new_n649), .ZN(new_n655));
  INV_X1    g454(.A(new_n584), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n652), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n651), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(G134gat), .B(G162gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AND4_X1   g462(.A1(new_n657), .A2(new_n658), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n658), .A2(new_n663), .B1(new_n660), .B2(new_n657), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n645), .A3(new_n639), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n644), .A2(new_n646), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n611), .A2(new_n613), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n612), .B1(new_n618), .B2(KEYINPUT97), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT101), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n614), .B(new_n619), .C1(new_n647), .C2(new_n649), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n671), .A2(new_n674), .A3(new_n672), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n650), .A2(new_n676), .A3(KEYINPUT10), .A4(new_n620), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n671), .A2(new_n674), .ZN(new_n681));
  INV_X1    g480(.A(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n680), .A2(new_n683), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n635), .A2(new_n666), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n608), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n523), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n538), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n575), .B2(new_n698), .ZN(new_n701));
  MUX2_X1   g500(.A(new_n700), .B(new_n701), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g501(.A(new_n498), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n695), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n535), .A2(G15gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n695), .B2(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n254), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n695), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NOR3_X1   g509(.A1(new_n635), .A2(new_n666), .A3(new_n691), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n608), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n517), .A3(new_n552), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n691), .B(KEYINPUT102), .Z(new_n716));
  NOR3_X1   g515(.A1(new_n635), .A2(new_n607), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n541), .B2(new_n666), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n530), .A2(new_n462), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n534), .A2(new_n540), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n666), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT44), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n718), .B1(new_n720), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n517), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n553), .B1(new_n729), .B2(KEYINPUT104), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n715), .B1(new_n730), .B2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n558), .A3(new_n437), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n558), .B1(new_n728), .B2(new_n437), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n728), .A2(new_n498), .ZN(new_n738));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n713), .A2(new_n739), .A3(new_n490), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  OAI221_X1 g543(.A(new_n741), .B1(new_n737), .B2(KEYINPUT47), .C1(new_n738), .C2(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1330gat));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n254), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n712), .A2(KEYINPUT106), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n707), .A2(G50gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n712), .B2(KEYINPUT106), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT48), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n747), .A2(G50gat), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n753), .A2(new_n755), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n752), .A2(new_n756), .B1(new_n759), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g559(.A(new_n635), .ZN(new_n761));
  INV_X1    g560(.A(new_n716), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n606), .A4(new_n724), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n723), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n523), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g565(.A(new_n764), .B(KEYINPUT108), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n538), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n498), .A2(G71gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n764), .A2(new_n535), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n767), .A2(new_n773), .B1(G71gat), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g575(.A1(new_n767), .A2(new_n707), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT109), .B(G78gat), .Z(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1335gat));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n541), .B2(new_n666), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n723), .A2(KEYINPUT110), .A3(new_n724), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n635), .A2(new_n606), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n783), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n666), .B1(new_n721), .B2(new_n722), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n637), .A3(new_n517), .A4(new_n691), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n720), .A2(new_n727), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n787), .A2(new_n692), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n523), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1336gat));
  INV_X1    g596(.A(new_n794), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n720), .B2(new_n727), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n638), .B1(new_n799), .B2(new_n437), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n762), .A2(new_n538), .A3(G92gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT52), .Z(G1337gat));
  NOR3_X1   g602(.A1(new_n535), .A2(G99gat), .A3(new_n692), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G99gat), .B1(new_n795), .B2(new_n703), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1338gat));
  NOR3_X1   g606(.A1(new_n762), .A2(new_n707), .A3(G106gat), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n786), .B2(new_n790), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(G106gat), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n799), .B2(new_n254), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n810), .A2(KEYINPUT112), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  AND4_X1   g615(.A1(KEYINPUT51), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n789), .B2(new_n781), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n808), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n795), .B2(new_n707), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n812), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n810), .B2(new_n814), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n816), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT53), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  NAND4_X1  g626(.A1(new_n635), .A2(new_n607), .A3(new_n666), .A4(new_n692), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n673), .A2(new_n675), .A3(new_n677), .A4(new_n682), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n680), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n678), .A2(new_n833), .A3(new_n679), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n688), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n829), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n688), .A4(new_n834), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n690), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n595), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n593), .A2(new_n588), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n586), .B1(new_n585), .B2(new_n588), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n586), .C1(new_n585), .C2(new_n588), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n601), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n605), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n666), .A2(new_n838), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n605), .A3(new_n691), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n607), .B2(new_n838), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n666), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n828), .B1(new_n850), .B2(new_n635), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n523), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n532), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n538), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n256), .A3(new_n606), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n437), .A2(new_n523), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n536), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n607), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT114), .Z(G1340gat));
  NOR3_X1   g661(.A1(new_n859), .A2(new_n258), .A3(new_n762), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n855), .A2(new_n691), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n258), .ZN(G1341gat));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n266), .A3(new_n635), .ZN(new_n866));
  OAI21_X1  g665(.A(G127gat), .B1(new_n859), .B2(new_n761), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT115), .Z(G1342gat));
  NOR2_X1   g668(.A1(new_n437), .A2(new_n666), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n264), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n859), .B2(new_n666), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  NOR2_X1   g674(.A1(new_n498), .A2(new_n707), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(G141gat), .A3(new_n607), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT58), .B1(new_n879), .B2(KEYINPUT122), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n851), .B2(new_n254), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n837), .A2(new_n690), .ZN(new_n883));
  INV_X1    g682(.A(new_n835), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT55), .B1(new_n884), .B2(new_n831), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT118), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n836), .A2(new_n887), .A3(new_n690), .A4(new_n837), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n606), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n845), .A2(new_n605), .A3(new_n891), .A4(new_n691), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n847), .B1(new_n893), .B2(new_n666), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n882), .B1(new_n894), .B2(new_n635), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n890), .A2(new_n892), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n724), .B1(new_n896), .B2(new_n889), .ZN(new_n897));
  OAI211_X1 g696(.A(KEYINPUT119), .B(new_n761), .C1(new_n897), .C2(new_n847), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n898), .A3(new_n828), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n254), .A2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n881), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n703), .A2(new_n857), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT116), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n607), .A3(new_n904), .ZN(new_n905));
  OAI221_X1 g704(.A(new_n880), .B1(KEYINPUT122), .B2(new_n879), .C1(new_n202), .C2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908));
  INV_X1    g707(.A(new_n904), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n761), .B1(new_n897), .B2(new_n847), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n910), .A2(new_n882), .B1(new_n607), .B2(new_n694), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n900), .B1(new_n911), .B2(new_n898), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n908), .B(new_n909), .C1(new_n912), .C2(new_n881), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n902), .B2(new_n904), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n606), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G141gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n879), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n907), .B1(new_n917), .B2(KEYINPUT58), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n878), .B1(new_n915), .B2(G141gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n906), .B1(new_n918), .B2(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(new_n877), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n204), .A3(new_n691), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n707), .B1(new_n910), .B2(new_n828), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .B1(new_n852), .B2(new_n900), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(new_n691), .A3(new_n909), .ZN(new_n927));
  NAND2_X1  g726(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n914), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n204), .B1(new_n930), .B2(new_n691), .ZN(new_n931));
  OAI221_X1 g730(.A(new_n924), .B1(new_n927), .B2(new_n928), .C1(new_n931), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g731(.A(G155gat), .B1(new_n929), .B2(new_n761), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n208), .A3(new_n635), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  NAND4_X1  g734(.A1(new_n853), .A2(new_n209), .A3(new_n870), .A4(new_n876), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n929), .B2(new_n666), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G162gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n929), .A2(KEYINPUT123), .A3(new_n666), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1347gat));
  NOR3_X1   g739(.A1(new_n852), .A2(new_n517), .A3(new_n538), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(new_n532), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n606), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n536), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n341), .A3(new_n607), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n943), .A2(new_n945), .ZN(G1348gat));
  AOI21_X1  g745(.A(G176gat), .B1(new_n942), .B2(new_n691), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n944), .A2(new_n342), .A3(new_n762), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n942), .A2(new_n388), .A3(new_n635), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n355), .A2(new_n356), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n944), .B2(new_n761), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n944), .B2(new_n666), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n331), .A3(new_n724), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n498), .A2(new_n517), .A3(new_n538), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT126), .Z(new_n961));
  NAND2_X1  g760(.A1(new_n926), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n607), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n851), .A2(new_n254), .A3(new_n960), .ZN(new_n964));
  INV_X1    g763(.A(G197gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(new_n606), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(G1352gat));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n969), .A3(new_n691), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n962), .B2(new_n762), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1353gat));
  NAND3_X1  g772(.A1(new_n964), .A2(new_n220), .A3(new_n635), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n926), .A2(new_n635), .A3(new_n961), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  AND2_X1   g777(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n724), .B1(new_n962), .B2(KEYINPUT127), .ZN(new_n980));
  OAI21_X1  g779(.A(G218gat), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n221), .A3(new_n724), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


