//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT70), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n460), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n466), .B2(new_n468), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n460), .A2(G138), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n463), .A2(new_n469), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n460), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n460), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n473), .A2(KEYINPUT71), .A3(G126), .A4(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n493), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT74), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n507), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n508), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n506), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT6), .B(G651), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(G50), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT75), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(G543), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(G543), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n506), .A2(new_n511), .A3(new_n515), .A4(new_n527), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n535), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n537), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n531), .A2(new_n533), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n516), .A2(G64), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n518), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n534), .A2(G43), .B1(G81), .B2(new_n537), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n518), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(KEYINPUT78), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND3_X1  g138(.A1(new_n529), .A2(KEYINPUT9), .A3(G53), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n532), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n506), .A2(new_n511), .A3(new_n515), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n537), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n518), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n537), .A2(G87), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n529), .A2(G49), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n536), .A2(new_n586), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n588), .B2(new_n580), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  NAND4_X1  g166(.A1(new_n506), .A2(new_n511), .A3(G86), .A4(new_n515), .ZN(new_n592));
  NAND2_X1  g167(.A1(G48), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n527), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n506), .A2(new_n511), .A3(G61), .A4(new_n515), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT81), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n537), .A2(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n546), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n516), .A2(G60), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n518), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(new_n518), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G54), .B2(new_n534), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n537), .A2(G92), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT10), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G868), .ZN(G321));
  XOR2_X1   g193(.A(G321), .B(KEYINPUT82), .Z(G284));
  MUX2_X1   g194(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n617), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND4_X1   g202(.A1(G2104), .A2(new_n463), .A3(new_n469), .A4(new_n460), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT12), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n482), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n479), .A2(KEYINPUT84), .A3(G135), .ZN(new_n640));
  AOI21_X1  g215(.A(KEYINPUT84), .B1(new_n479), .B2(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n637), .B1(new_n638), .B2(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n633), .B2(new_n634), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n636), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT14), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(new_n660), .A3(G14), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(KEYINPUT17), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n665), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n665), .B1(new_n662), .B2(new_n663), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n668), .B2(new_n662), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  OAI221_X1 g249(.A(new_n667), .B1(new_n668), .B2(new_n669), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n634), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G168), .A2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT94), .Z(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G16), .B2(G21), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1966), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G5), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G171), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G33), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n708));
  NAND2_X1  g283(.A1(G103), .A2(G2104), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n479), .A2(G139), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n463), .A2(new_n469), .A3(G127), .ZN(new_n713));
  NAND2_X1  g288(.A1(G115), .A2(G2104), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n460), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n707), .B1(new_n718), .B2(new_n706), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2072), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n705), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n706), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n706), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  INV_X1    g301(.A(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n726), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G160), .B2(new_n706), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n733));
  INV_X1    g308(.A(G141), .ZN(new_n734));
  INV_X1    g309(.A(G129), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n733), .B1(new_n478), .B2(new_n734), .C1(new_n735), .C2(new_n481), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n706), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n706), .B2(G32), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n706), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  INV_X1    g322(.A(G104), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n748), .A2(new_n460), .A3(KEYINPUT90), .ZN(new_n749));
  AOI21_X1  g324(.A(KEYINPUT90), .B1(new_n748), .B2(new_n460), .ZN(new_n750));
  OAI221_X1 g325(.A(G2104), .B1(G116), .B2(new_n460), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G128), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n753), .A2(new_n481), .B1(new_n478), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n747), .B1(new_n757), .B2(new_n706), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n743), .A2(new_n744), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n745), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n706), .A2(G35), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT95), .Z(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n706), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT29), .B(G2090), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n642), .A2(new_n706), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n769), .A2(G28), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n706), .B1(new_n769), .B2(G28), .ZN(new_n771));
  AND2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n767), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n765), .A2(new_n766), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n775), .B(new_n776), .C1(G2084), .C2(new_n730), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n721), .A2(new_n732), .A3(new_n762), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n701), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n617), .B2(new_n701), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1348), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n701), .A2(G20), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT23), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n701), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n558), .B2(new_n701), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1341), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n700), .A2(new_n778), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n706), .A2(G25), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n479), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n482), .A2(G119), .ZN(new_n795));
  OR2_X1    g370(.A1(G95), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT86), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(new_n706), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XOR2_X1   g377(.A(new_n801), .B(new_n802), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n608), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G16), .B2(G24), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n689), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n689), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n803), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT87), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n811), .B(KEYINPUT87), .ZN(new_n815));
  INV_X1    g390(.A(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n814), .A2(new_n817), .A3(KEYINPUT88), .ZN(new_n821));
  NOR2_X1   g396(.A1(G166), .A2(new_n701), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n701), .B2(G22), .ZN(new_n823));
  INV_X1    g398(.A(G1971), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n701), .A2(G23), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n588), .A2(new_n580), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n701), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT33), .B(G1976), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n823), .A2(new_n824), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n820), .A2(new_n821), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n810), .B1(new_n835), .B2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT89), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n820), .A2(new_n834), .A3(new_n838), .A4(new_n821), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n836), .B2(new_n839), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n792), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(new_n839), .A3(new_n809), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT89), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .A3(new_n840), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n791), .B1(new_n843), .B2(new_n847), .ZN(G311));
  INV_X1    g423(.A(new_n791), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n846), .A2(KEYINPUT36), .A3(new_n840), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT36), .B1(new_n846), .B2(new_n840), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(G150));
  NAND2_X1  g427(.A1(new_n537), .A2(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n516), .A2(G67), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n518), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n853), .B1(new_n546), .B2(new_n854), .C1(new_n857), .C2(KEYINPUT96), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(KEYINPUT96), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT98), .B(G860), .Z(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n558), .A2(new_n860), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n556), .A2(new_n557), .B1(new_n859), .B2(new_n858), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n616), .A2(new_n622), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n867), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n870), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT99), .B1(new_n870), .B2(new_n871), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n861), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n863), .B1(new_n874), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n642), .B(G160), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n479), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n482), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(G106), .A2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n632), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n798), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n891), .A2(KEYINPUT101), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT101), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n501), .B1(new_n493), .B2(KEYINPUT100), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n897));
  AOI211_X1 g472(.A(new_n897), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n757), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n741), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(new_n718), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n718), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n882), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n892), .A3(new_n891), .ZN(new_n909));
  INV_X1    g484(.A(new_n882), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n893), .A2(new_n894), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n904), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n882), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n911), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g497(.A(new_n866), .B(new_n624), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n617), .A2(G299), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n616), .A2(new_n574), .A3(new_n569), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n926), .B2(new_n923), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n608), .B(G305), .ZN(new_n933));
  XOR2_X1   g508(.A(G166), .B(new_n827), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n932), .A2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G868), .B2(new_n860), .ZN(G295));
  OAI21_X1  g515(.A(new_n939), .B1(G868), .B2(new_n860), .ZN(G331));
  XOR2_X1   g516(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n942));
  XNOR2_X1  g517(.A(new_n935), .B(KEYINPUT105), .ZN(new_n943));
  NAND2_X1  g518(.A1(G286), .A2(G301), .ZN(new_n944));
  NAND2_X1  g519(.A1(G168), .A2(G171), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n866), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n864), .A2(new_n865), .A3(new_n944), .A4(new_n945), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n866), .A2(new_n950), .A3(new_n946), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n926), .B(new_n927), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n949), .A2(new_n926), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n947), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n943), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n948), .A3(new_n951), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n960), .A3(new_n935), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n912), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n957), .A2(new_n962), .A3(KEYINPUT43), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n866), .A2(new_n950), .A3(new_n946), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n950), .B1(new_n866), .B2(new_n946), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n967), .A2(new_n955), .B1(new_n953), .B2(new_n959), .ZN(new_n968));
  AOI21_X1  g543(.A(G37), .B1(new_n968), .B2(new_n935), .ZN(new_n969));
  INV_X1    g544(.A(new_n943), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n958), .A2(new_n960), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n964), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n942), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n964), .A3(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n957), .B2(new_n962), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n472), .A2(new_n983), .A3(new_n476), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n896), .B2(new_n898), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n980), .B1(new_n988), .B2(G1966), .ZN(new_n989));
  INV_X1    g564(.A(G1966), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n491), .A2(new_n492), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n897), .B1(new_n991), .B2(new_n489), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n493), .A2(KEYINPUT100), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n501), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n994), .B2(new_n981), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT112), .B(new_n990), .C1(new_n995), .C2(new_n985), .ZN(new_n996));
  INV_X1    g571(.A(new_n476), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n470), .A2(new_n471), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(G40), .B(new_n997), .C1(new_n999), .C2(new_n460), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n502), .A2(new_n981), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2084), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n981), .C1(new_n896), .C2(new_n898), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n989), .A2(new_n996), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n979), .B1(new_n1007), .B2(G286), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n989), .A2(G168), .A3(new_n996), .A4(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n979), .B1(new_n1009), .B2(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT121), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(KEYINPUT51), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(new_n1015), .C1(new_n1010), .C2(new_n1008), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(KEYINPUT62), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT124), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1013), .A2(KEYINPUT124), .A3(new_n1016), .A4(KEYINPUT62), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT62), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1016), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n990), .B1(new_n995), .B2(new_n985), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n980), .ZN(new_n1025));
  AOI21_X1  g600(.A(G168), .B1(new_n1025), .B2(new_n996), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1009), .C1(new_n1026), .C2(new_n979), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1015), .B1(new_n1027), .B2(new_n1014), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1021), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n519), .B2(new_n523), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1030), .B(KEYINPUT55), .Z(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1001), .A2(new_n1033), .A3(new_n986), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT45), .B(new_n981), .C1(new_n896), .C2(new_n898), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n493), .B2(new_n501), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT110), .B1(new_n1036), .B2(KEYINPUT45), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n984), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n824), .ZN(new_n1039));
  INV_X1    g614(.A(G2090), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1002), .A2(new_n1040), .A3(new_n1005), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1032), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1031), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n984), .B(new_n981), .C1(new_n896), .C2(new_n898), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n827), .A2(G1976), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n585), .A2(new_n1048), .A3(new_n589), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n694), .B1(new_n595), .B2(new_n600), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n520), .B1(new_n592), .B2(new_n593), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n518), .B1(new_n596), .B2(new_n598), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1053), .A2(new_n1054), .A3(G1981), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1051), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n595), .A2(new_n600), .A3(new_n694), .ZN(new_n1057));
  OAI21_X1  g632(.A(G1981), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT49), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1045), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(G8), .A3(new_n1044), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1050), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1004), .B1(new_n994), .B2(new_n981), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n984), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT111), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1000), .B1(new_n1004), .B2(new_n1036), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1040), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1032), .B1(new_n1072), .B2(new_n1039), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1043), .B(new_n1064), .C1(new_n1073), .C2(new_n1031), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1038), .B2(G2078), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n988), .A2(KEYINPUT53), .A3(new_n724), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n704), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1019), .A2(new_n1020), .A3(new_n1029), .A4(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1044), .A2(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(new_n616), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(KEYINPUT60), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1044), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT120), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1038), .A2(G1996), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n558), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n558), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT56), .B(G2072), .Z(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1038), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n785), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(new_n785), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n574), .A2(new_n567), .A3(new_n564), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(G299), .C2(new_n1109), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1107), .A2(new_n1113), .A3(KEYINPUT61), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT61), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1089), .B(new_n1098), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1086), .A2(new_n616), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT119), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1074), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1080), .B2(G301), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT106), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT45), .B1(new_n987), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n981), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR4_X1   g703(.A1(new_n476), .A2(new_n1075), .A3(new_n983), .A4(G2078), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n998), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(G2105), .B1(new_n999), .B2(KEYINPUT122), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1035), .B(new_n1129), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1076), .B(new_n1079), .C1(new_n1128), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G171), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(KEYINPUT123), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1124), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1081), .B(new_n1123), .C1(G171), .C2(new_n1134), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1122), .A2(new_n1013), .A3(new_n1016), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1042), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1031), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT114), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G286), .A2(new_n1032), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1007), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1063), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1042), .B1(new_n1031), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(G2090), .B1(new_n1102), .B2(KEYINPUT111), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1153), .A2(new_n1071), .B1(new_n824), .B2(new_n1038), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1143), .B1(new_n1154), .B2(new_n1032), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1063), .B1(new_n1031), .B2(new_n1042), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1146), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1155), .A2(new_n1156), .A3(new_n1146), .A4(KEYINPUT113), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1045), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n1048), .A3(new_n590), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1164), .B2(new_n1057), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1043), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1064), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT115), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1146), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1158), .B1(new_n1074), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1171), .A2(new_n1147), .A3(new_n1160), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1151), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT115), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n1174), .A3(new_n1167), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1083), .A2(new_n1141), .A3(new_n1169), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1128), .A2(new_n984), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n608), .A2(new_n689), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT107), .Z(new_n1182));
  INV_X1    g757(.A(G1996), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1178), .A2(KEYINPUT108), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT108), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1177), .B2(G1996), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n756), .B(new_n759), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1183), .B2(new_n741), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1187), .A2(new_n741), .B1(new_n1178), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n798), .B(new_n802), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n1178), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1182), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT109), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1176), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1187), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1184), .A2(KEYINPUT46), .A3(new_n1186), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1177), .B1(new_n741), .B2(new_n1188), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(KEYINPUT126), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1199), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1203), .A2(KEYINPUT47), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1190), .A2(new_n800), .A3(new_n802), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(G2067), .B2(new_n756), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1178), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1190), .A2(new_n1192), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1206), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT47), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1195), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g791(.A1(new_n963), .A2(new_n973), .ZN(new_n1218));
  INV_X1    g792(.A(new_n458), .ZN(new_n1219));
  NOR2_X1   g793(.A1(G227), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g794(.A(new_n1220), .B(KEYINPUT127), .ZN(new_n1221));
  NOR3_X1   g795(.A1(new_n1221), .A2(G401), .A3(G229), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n921), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n1218), .A2(new_n1223), .ZN(G308));
  OAI211_X1 g798(.A(new_n921), .B(new_n1222), .C1(new_n963), .C2(new_n973), .ZN(G225));
endmodule


