//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  OR2_X1    g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G57gat), .A2(G64gat), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n204), .C1(new_n207), .C2(KEYINPUT9), .ZN(new_n208));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT96), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(new_n209), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT97), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(G231gat), .A2(G233gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(G231gat), .B(G233gat), .C1(new_n219), .C2(KEYINPUT21), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(KEYINPUT20), .Z(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n225), .A2(new_n227), .ZN(new_n229));
  XOR2_X1   g028(.A(G183gat), .B(G211gat), .Z(new_n230));
  OR3_X1    g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G15gat), .B(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT92), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n232), .A2(new_n233), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n235), .A2(G1gat), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G1gat), .ZN(new_n239));
  XOR2_X1   g038(.A(G15gat), .B(G22gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT92), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n241), .B2(new_n234), .ZN(new_n242));
  OAI21_X1  g041(.A(G8gat), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  OAI22_X1  g042(.A1(new_n235), .A2(new_n236), .B1(new_n238), .B2(G1gat), .ZN(new_n244));
  INV_X1    g043(.A(G8gat), .ZN(new_n245));
  INV_X1    g044(.A(G1gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n246), .A3(new_n234), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n220), .B2(new_n221), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  OAI21_X1  g052(.A(new_n230), .B1(new_n228), .B2(new_n229), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n231), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n231), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT15), .ZN(new_n259));
  INV_X1    g058(.A(G50gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G43gat), .ZN(new_n261));
  INV_X1    g060(.A(G43gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G50gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT88), .ZN(new_n267));
  NAND2_X1  g066(.A1(G29gat), .A2(G36gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR3_X1   g069(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n271), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT91), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n276), .B2(KEYINPUT91), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n277), .A2(new_n278), .B1(new_n266), .B2(new_n267), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT90), .B(G50gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n261), .B1(new_n280), .B2(G43gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n281), .A2(new_n259), .B1(G29gat), .B2(G36gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT17), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT94), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n273), .A2(new_n274), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n273), .A2(new_n274), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(new_n288), .B1(new_n282), .B2(new_n279), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT17), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n285), .ZN(new_n293));
  NAND2_X1  g092(.A1(G85gat), .A2(G92gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT7), .ZN(new_n295));
  NOR2_X1   g094(.A1(G85gat), .A2(G92gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G99gat), .A2(G106gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(KEYINPUT8), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G99gat), .B(G106gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n292), .A2(new_n293), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n301), .ZN(new_n303));
  AND2_X1   g102(.A1(G232gat), .A2(G233gat), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n284), .A2(new_n303), .B1(KEYINPUT41), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G190gat), .B(G218gat), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n304), .A2(KEYINPUT41), .ZN(new_n312));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(new_n314), .A3(new_n310), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT100), .ZN(new_n323));
  INV_X1    g122(.A(G230gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n301), .A2(new_n213), .A3(new_n218), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n299), .A2(KEYINPUT99), .ZN(new_n329));
  INV_X1    g128(.A(new_n300), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n299), .A2(KEYINPUT99), .A3(new_n300), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n331), .B(new_n332), .C1(new_n212), .C2(new_n211), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n303), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n327), .B2(new_n333), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n323), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n339), .A2(KEYINPUT101), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(KEYINPUT101), .ZN(new_n341));
  INV_X1    g140(.A(new_n336), .ZN(new_n342));
  INV_X1    g141(.A(new_n338), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n322), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n258), .A2(new_n319), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347));
  NAND2_X1  g146(.A1(G211gat), .A2(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(G211gat), .ZN(new_n349));
  INV_X1    g148(.A(G218gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(G197gat), .A2(G204gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n348), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n348), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n348), .A2(new_n355), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G226gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n325), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT23), .ZN(new_n370));
  INV_X1    g169(.A(G169gat), .ZN(new_n371));
  INV_X1    g170(.A(G176gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  NOR2_X1   g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT23), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n368), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n366), .A2(new_n380), .A3(new_n367), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n366), .B2(new_n367), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n372), .ZN(new_n385));
  NAND2_X1  g184(.A1(KEYINPUT67), .A2(G176gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(KEYINPUT23), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n371), .A2(KEYINPUT66), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT66), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G169gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n374), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT68), .B(new_n374), .C1(new_n387), .C2(new_n391), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n383), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n379), .B1(new_n396), .B2(new_n375), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT70), .B(KEYINPUT26), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT71), .B1(new_n398), .B2(new_n373), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT26), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n376), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n369), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(KEYINPUT26), .B2(new_n373), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G183gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT27), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G183gat), .ZN(new_n411));
  INV_X1    g210(.A(G190gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT28), .A4(new_n412), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT69), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n418), .A3(new_n414), .ZN(new_n419));
  AND4_X1   g218(.A1(new_n365), .A2(new_n407), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n363), .B1(new_n397), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT76), .B(new_n363), .C1(new_n397), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n397), .B2(new_n420), .ZN(new_n427));
  INV_X1    g226(.A(new_n363), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n361), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n361), .A3(new_n421), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT77), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT77), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n423), .A2(new_n424), .B1(new_n428), .B2(new_n427), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n434), .B(new_n431), .C1(new_n435), .C2(new_n361), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n433), .A2(KEYINPUT78), .A3(new_n436), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT31), .B(G50gat), .ZN(new_n446));
  XOR2_X1   g245(.A(G141gat), .B(G148gat), .Z(new_n447));
  INV_X1    g246(.A(G155gat), .ZN(new_n448));
  INV_X1    g247(.A(G162gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(KEYINPUT2), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G141gat), .B(G148gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n451), .B(new_n450), .C1(new_n455), .C2(KEYINPUT2), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n356), .B2(new_n360), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(KEYINPUT82), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n462), .B(KEYINPUT29), .C1(new_n356), .C2(new_n360), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n458), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(new_n456), .A3(new_n459), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n361), .B1(new_n465), .B2(new_n426), .ZN(new_n466));
  NAND2_X1  g265(.A1(G228gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  INV_X1    g270(.A(new_n360), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n357), .B1(new_n359), .B2(new_n358), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n426), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n457), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n470), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n471), .B1(new_n470), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n446), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n459), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n474), .B2(new_n462), .ZN(new_n482));
  INV_X1    g281(.A(new_n463), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n457), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n466), .A2(new_n468), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n477), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n477), .ZN(new_n488));
  INV_X1    g287(.A(new_n446), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(G22gat), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n480), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n480), .B2(new_n490), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n396), .A2(new_n375), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n420), .B1(new_n496), .B2(new_n378), .ZN(new_n497));
  XNOR2_X1  g296(.A(G113gat), .B(G120gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT1), .ZN(new_n501));
  XNOR2_X1  g300(.A(G127gat), .B(G134gat), .ZN(new_n502));
  INV_X1    g301(.A(G113gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n502), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(KEYINPUT1), .B2(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT64), .Z(new_n511));
  AND3_X1   g310(.A1(new_n502), .A2(new_n501), .A3(new_n504), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n498), .A2(KEYINPUT1), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n512), .A2(new_n500), .B1(new_n513), .B2(new_n506), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n397), .B2(new_n420), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G43gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT73), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G71gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(G99gat), .Z(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n523), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT32), .B(new_n516), .C1(new_n525), .C2(new_n518), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n511), .A2(KEYINPUT34), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n509), .B2(new_n515), .ZN(new_n528));
  INV_X1    g327(.A(new_n515), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n397), .A2(new_n420), .A3(new_n514), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n510), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n531), .B2(KEYINPUT34), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n524), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n524), .B2(new_n526), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n495), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n431), .B(new_n439), .C1(new_n435), .C2(new_n361), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT30), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT81), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n505), .A2(new_n456), .A3(new_n454), .A4(new_n507), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT4), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT4), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n541), .A4(new_n457), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n508), .B(new_n465), .C1(new_n457), .C2(new_n475), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT5), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G225gat), .A2(G233gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n514), .A2(new_n457), .A3(new_n543), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n539), .A2(new_n541), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT5), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n508), .B(new_n457), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n548), .A2(new_n553), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n547), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G1gat), .B(G29gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT0), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G85gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  AOI21_X1  g360(.A(KEYINPUT6), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n554), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n561), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(KEYINPUT6), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n445), .A2(new_n535), .A3(new_n537), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT35), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n575));
  INV_X1    g374(.A(new_n495), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n524), .A2(new_n526), .ZN(new_n578));
  INV_X1    g377(.A(new_n532), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n524), .A2(new_n526), .A3(new_n532), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n581), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n534), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n576), .B(new_n577), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n445), .A2(new_n537), .A3(new_n570), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n574), .A2(new_n575), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n433), .A2(KEYINPUT37), .A3(new_n436), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n591));
  OAI211_X1 g390(.A(new_n431), .B(new_n591), .C1(new_n435), .C2(new_n361), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n592), .A2(new_n440), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT38), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n568), .A2(new_n536), .A3(new_n569), .ZN(new_n596));
  INV_X1    g395(.A(new_n361), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n429), .A2(new_n597), .A3(new_n421), .ZN(new_n598));
  OAI211_X1 g397(.A(KEYINPUT37), .B(new_n598), .C1(new_n435), .C2(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n596), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n495), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n536), .B(KEYINPUT30), .Z(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n443), .B2(new_n444), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n552), .A2(new_n549), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n555), .A2(new_n548), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(KEYINPUT39), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n561), .C1(KEYINPUT39), .C2(new_n606), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT40), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n567), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n603), .B(KEYINPUT85), .C1(new_n605), .C2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT85), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n445), .B2(new_n537), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n600), .B1(new_n590), .B2(new_n593), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n592), .A2(new_n599), .A3(new_n600), .A4(new_n440), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n536), .A3(new_n568), .A4(new_n569), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n576), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n613), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n580), .A2(KEYINPUT36), .A3(new_n582), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n534), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n587), .A2(new_n495), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n612), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n589), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT93), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n237), .A2(new_n242), .A3(G8gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n245), .B1(new_n244), .B2(new_n247), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n243), .A2(KEYINPUT93), .A3(new_n248), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n284), .A2(KEYINPUT94), .A3(new_n285), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n290), .B1(new_n289), .B2(KEYINPUT17), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n639), .B(new_n293), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G229gat), .A2(G233gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n250), .A2(new_n289), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n284), .B(new_n249), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n643), .B(KEYINPUT13), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n637), .A2(new_n638), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n289), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n644), .B1(new_n292), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT18), .B1(new_n654), .B2(new_n643), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n633), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n633), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n646), .A3(new_n649), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n347), .B1(new_n627), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n656), .A2(new_n661), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT95), .B(new_n664), .C1(new_n589), .C2(new_n626), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n346), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n570), .B(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  INV_X1    g469(.A(new_n605), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(new_n346), .C1(new_n663), .C2(new_n665), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(G8gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT42), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n624), .A2(new_n620), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n666), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n583), .A2(new_n585), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n666), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n495), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n345), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n258), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n318), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n627), .A2(new_n662), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT95), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n627), .A2(new_n347), .A3(new_n662), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n668), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(G29gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n627), .A2(new_n319), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n627), .A2(KEYINPUT44), .A3(new_n319), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n664), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n697), .A2(KEYINPUT45), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n698), .B1(new_n706), .B2(new_n707), .ZN(G1328gat));
  INV_X1    g507(.A(G36gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n709), .A3(new_n671), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n705), .B2(new_n605), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(KEYINPUT46), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(new_n690), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n663), .B2(new_n665), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n262), .B1(new_n716), .B2(new_n681), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n679), .A2(new_n262), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n704), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n495), .A2(new_n280), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(KEYINPUT105), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(KEYINPUT105), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n694), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n701), .A2(new_n495), .A3(new_n702), .A4(new_n704), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n280), .A2(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n729), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1331gat));
  NOR4_X1   g535(.A1(new_n258), .A2(new_n319), .A3(new_n662), .A4(new_n687), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n627), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n668), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n739), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n605), .B(KEYINPUT108), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n739), .B(KEYINPUT107), .ZN(new_n752));
  INV_X1    g551(.A(new_n679), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n205), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n739), .A2(G71gat), .A3(new_n681), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G71gat), .B1(new_n744), .B2(new_n679), .ZN(new_n757));
  INV_X1    g556(.A(new_n755), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(KEYINPUT50), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n752), .A2(new_n495), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n695), .A2(G85gat), .A3(new_n687), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n257), .A2(new_n662), .ZN(new_n764));
  INV_X1    g563(.A(new_n575), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT86), .B1(new_n571), .B2(KEYINPUT35), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n586), .A2(new_n587), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n612), .A2(new_n619), .A3(new_n625), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n319), .B(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n627), .A2(KEYINPUT51), .A3(new_n319), .A4(new_n764), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(KEYINPUT110), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n775), .A3(new_n771), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT111), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n763), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n257), .A2(new_n662), .A3(new_n687), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n701), .A2(new_n668), .A3(new_n702), .A4(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(G85gat), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n785), .ZN(G1336gat));
  INV_X1    g585(.A(new_n745), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n701), .A2(new_n702), .A3(new_n787), .A4(new_n780), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n745), .A2(G92gat), .A3(new_n687), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n774), .A2(new_n776), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n701), .A2(new_n671), .A3(new_n702), .A4(new_n780), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n773), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(G92gat), .B1(new_n795), .B2(new_n792), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n793), .B1(new_n796), .B2(new_n790), .ZN(G1337gat));
  NOR3_X1   g596(.A1(new_n681), .A2(new_n687), .A3(G99gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n777), .B2(new_n778), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n703), .A2(new_n753), .A3(new_n780), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1338gat));
  NAND4_X1  g601(.A1(new_n701), .A2(new_n495), .A3(new_n702), .A4(new_n780), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n576), .A2(G106gat), .A3(new_n687), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n774), .A2(new_n776), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n803), .A2(G106gat), .B1(new_n795), .B2(new_n807), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n806), .A2(new_n808), .B1(new_n809), .B2(new_n805), .ZN(G1339gat));
  NAND2_X1  g609(.A1(new_n346), .A2(new_n664), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n334), .A2(new_n335), .A3(new_n326), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT112), .A4(new_n326), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n342), .A3(KEYINPUT54), .A4(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n322), .B1(new_n336), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n344), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT113), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n822), .A3(new_n344), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(new_n816), .B2(new_n818), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n654), .A2(new_n643), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n647), .A2(new_n648), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n632), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n661), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n826), .A2(new_n318), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n661), .A2(new_n345), .A3(new_n829), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n661), .A2(new_n829), .A3(KEYINPUT114), .A4(new_n345), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n834), .B(new_n835), .C1(new_n826), .C2(new_n664), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n831), .B1(new_n836), .B2(new_n318), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n811), .B1(new_n837), .B2(new_n257), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n668), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n745), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n681), .A2(new_n495), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n662), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(G113gat), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n842), .B2(G113gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n535), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n662), .A2(new_n503), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n845), .A2(new_n846), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  OR3_X1    g648(.A1(new_n847), .A2(G120gat), .A3(new_n687), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n840), .A2(new_n841), .A3(new_n345), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n851), .B2(G120gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n841), .A3(new_n257), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G127gat), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n258), .A2(G127gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n847), .B2(new_n858), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n671), .A2(new_n318), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n839), .A2(new_n860), .A3(new_n535), .A4(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT56), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n841), .A3(new_n319), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(G134gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n864), .B2(G134gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n753), .A2(new_n576), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n839), .A2(new_n745), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n664), .A2(G141gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n838), .A2(new_n874), .A3(new_n495), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n745), .A2(new_n679), .A3(new_n668), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n820), .B2(new_n824), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n825), .A2(KEYINPUT118), .A3(new_n344), .A4(new_n819), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n662), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n319), .B1(new_n880), .B2(new_n832), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n258), .B1(new_n881), .B2(new_n831), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n576), .B1(new_n882), .B2(new_n811), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n876), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n662), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n873), .B1(new_n886), .B2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n873), .B2(KEYINPUT119), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(G1344gat));
  OR3_X1    g688(.A1(new_n871), .A2(G148gat), .A3(new_n687), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n838), .A2(new_n495), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n883), .A2(new_n874), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n345), .A3(new_n876), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(G148gat), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n885), .B2(new_n345), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n890), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n890), .B(new_n901), .C1(new_n896), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1345gat));
  NOR2_X1   g702(.A1(new_n871), .A2(new_n258), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g704(.A(G155gat), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n258), .A2(new_n448), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(new_n885), .B2(new_n907), .ZN(G1346gat));
  NAND4_X1  g707(.A1(new_n839), .A2(new_n449), .A3(new_n861), .A4(new_n870), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n875), .A2(new_n884), .A3(new_n318), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n449), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n745), .A2(new_n668), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n838), .A2(new_n912), .A3(new_n535), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(new_n662), .A3(new_n388), .A4(new_n390), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n671), .A2(new_n695), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT122), .B1(new_n915), .B2(new_n681), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n681), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n576), .A2(new_n838), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n662), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n914), .B1(new_n371), .B2(new_n919), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n913), .B2(new_n345), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n687), .B1(new_n385), .B2(new_n386), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n918), .B2(new_n922), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n257), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G183gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n913), .A2(new_n409), .A3(new_n411), .A4(new_n257), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n932), .B(new_n925), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  AOI21_X1  g733(.A(new_n412), .B1(new_n918), .B2(new_n319), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT61), .Z(new_n936));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n412), .A3(new_n319), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1351gat));
  AND3_X1   g737(.A1(new_n838), .A2(new_n912), .A3(new_n870), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n662), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n893), .A2(new_n894), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n671), .A2(new_n679), .A3(new_n695), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n942), .A2(new_n664), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n944), .B2(new_n940), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(new_n941), .C1(new_n944), .C2(new_n940), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(G204gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n939), .A2(new_n950), .A3(new_n345), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(KEYINPUT62), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(KEYINPUT125), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT62), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n942), .A2(new_n687), .A3(new_n943), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n956), .C1(new_n950), .C2(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n874), .B1(new_n838), .B2(new_n495), .ZN(new_n961));
  AOI211_X1 g760(.A(KEYINPUT57), .B(new_n576), .C1(new_n882), .C2(new_n811), .ZN(new_n962));
  NOR4_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n258), .A4(new_n943), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n349), .B1(KEYINPUT126), .B2(new_n959), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n960), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n943), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n893), .A2(new_n257), .A3(new_n894), .A4(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n960), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n964), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n939), .A2(new_n349), .A3(new_n257), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n966), .A2(KEYINPUT127), .A3(new_n970), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n939), .A2(new_n350), .A3(new_n319), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n942), .A2(new_n318), .A3(new_n943), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n350), .ZN(G1355gat));
endmodule


