

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(KEYINPUT13), .ZN(n590) );
  OR2_X1 U555 ( .A1(n762), .A2(n761), .ZN(n520) );
  OR2_X1 U556 ( .A1(n764), .A2(n778), .ZN(n521) );
  XOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .Z(n522) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n694) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n719) );
  XNOR2_X1 U560 ( .A(n720), .B(n719), .ZN(n726) );
  XNOR2_X1 U561 ( .A(n746), .B(KEYINPUT32), .ZN(n770) );
  AND2_X1 U562 ( .A1(n1007), .A2(n521), .ZN(n765) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n795) );
  NOR2_X1 U564 ( .A1(n661), .A2(n539), .ZN(n647) );
  XNOR2_X1 U565 ( .A(n527), .B(KEYINPUT65), .ZN(n891) );
  NOR2_X1 U566 ( .A1(G651), .A2(n661), .ZN(n656) );
  INV_X1 U567 ( .A(G2104), .ZN(n523) );
  NOR2_X1 U568 ( .A1(G2105), .A2(n523), .ZN(n576) );
  BUF_X1 U569 ( .A(n576), .Z(n894) );
  NAND2_X1 U570 ( .A1(G102), .A2(n894), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n524), .Z(n895) );
  NAND2_X1 U573 ( .A1(G138), .A2(n895), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n523), .A2(G2105), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G126), .A2(n891), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT66), .B(n528), .Z(n781) );
  NAND2_X1 U579 ( .A1(G114), .A2(n781), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(G164) );
  XOR2_X1 U582 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n534) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U584 ( .A1(G89), .A2(n650), .ZN(n533) );
  XNOR2_X1 U585 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT72), .B(n535), .ZN(n537) );
  XNOR2_X1 U587 ( .A(KEYINPUT68), .B(n522), .ZN(n661) );
  INV_X1 U588 ( .A(G651), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n647), .A2(G76), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n538), .B(KEYINPUT5), .ZN(n545) );
  NOR2_X1 U592 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n540), .Z(n660) );
  NAND2_X1 U594 ( .A1(G63), .A2(n660), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G51), .A2(n656), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U599 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U601 ( .A(G2454), .B(G2446), .ZN(n556) );
  XOR2_X1 U602 ( .A(G2430), .B(KEYINPUT104), .Z(n548) );
  XNOR2_X1 U603 ( .A(G2451), .B(G2443), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n548), .B(n547), .ZN(n552) );
  XOR2_X1 U605 ( .A(G2427), .B(KEYINPUT103), .Z(n550) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U608 ( .A(n552), .B(n551), .Z(n554) );
  XNOR2_X1 U609 ( .A(G2435), .B(G2438), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U612 ( .A1(n557), .A2(G14), .ZN(G401) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G123), .A2(n891), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT18), .ZN(n565) );
  NAND2_X1 U616 ( .A1(G99), .A2(n894), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G135), .A2(n895), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n781), .A2(G111), .ZN(n561) );
  XOR2_X1 U620 ( .A(KEYINPUT76), .B(n561), .Z(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U623 ( .A(KEYINPUT77), .B(n566), .Z(n920) );
  XNOR2_X1 U624 ( .A(G2096), .B(n920), .ZN(n567) );
  OR2_X1 U625 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  NAND2_X1 U629 ( .A1(G64), .A2(n660), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(KEYINPUT69), .ZN(n575) );
  NAND2_X1 U631 ( .A1(G90), .A2(n650), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G77), .A2(n647), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n571), .B(KEYINPUT9), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G52), .A2(n656), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U638 ( .A1(n895), .A2(G137), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G101), .A2(n576), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n577), .Z(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G125), .A2(n891), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G113), .A2(n781), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n583), .A2(n582), .ZN(G160) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U647 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n837) );
  NAND2_X1 U649 ( .A1(n837), .A2(G567), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U651 ( .A1(G56), .A2(n660), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT14), .B(n586), .Z(n593) );
  NAND2_X1 U653 ( .A1(G68), .A2(n647), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n650), .A2(G81), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n591), .B(n590), .ZN(n592) );
  NOR2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n656), .A2(G43), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n994) );
  INV_X1 U661 ( .A(G860), .ZN(n617) );
  NOR2_X1 U662 ( .A1(n994), .A2(n617), .ZN(n596) );
  XOR2_X1 U663 ( .A(KEYINPUT70), .B(n596), .Z(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U666 ( .A1(n647), .A2(G79), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G92), .A2(n650), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G66), .A2(n660), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G54), .A2(n656), .ZN(n599) );
  XNOR2_X1 U671 ( .A(KEYINPUT71), .B(n599), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U674 ( .A(KEYINPUT15), .B(n604), .Z(n705) );
  INV_X1 U675 ( .A(G868), .ZN(n675) );
  NAND2_X1 U676 ( .A1(n705), .A2(n675), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G65), .A2(n660), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G53), .A2(n656), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G91), .A2(n650), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G78), .A2(n647), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n715) );
  INV_X1 U685 ( .A(n715), .ZN(G299) );
  XNOR2_X1 U686 ( .A(KEYINPUT74), .B(n675), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G286), .A2(n613), .ZN(n615) );
  NOR2_X1 U688 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U690 ( .A(KEYINPUT75), .B(n616), .Z(G297) );
  NAND2_X1 U691 ( .A1(n617), .A2(G559), .ZN(n618) );
  INV_X1 U692 ( .A(n705), .ZN(n993) );
  NAND2_X1 U693 ( .A1(n618), .A2(n993), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(G868), .A2(n994), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G868), .A2(n993), .ZN(n620) );
  NOR2_X1 U697 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G93), .A2(n650), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G67), .A2(n660), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G80), .A2(n647), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G55), .A2(n656), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n676) );
  XNOR2_X1 U706 ( .A(KEYINPUT78), .B(n994), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n993), .A2(G559), .ZN(n672) );
  XNOR2_X1 U708 ( .A(n629), .B(n672), .ZN(n630) );
  NOR2_X1 U709 ( .A1(G860), .A2(n630), .ZN(n631) );
  XOR2_X1 U710 ( .A(n676), .B(n631), .Z(G145) );
  NAND2_X1 U711 ( .A1(G86), .A2(n650), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G61), .A2(n660), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n647), .A2(G73), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n656), .A2(G48), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U719 ( .A1(G62), .A2(n660), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT80), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G75), .A2(n647), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G50), .A2(n656), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G88), .A2(n650), .ZN(n642) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n642), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(G303) );
  INV_X1 U728 ( .A(G303), .ZN(G166) );
  NAND2_X1 U729 ( .A1(G72), .A2(n647), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G47), .A2(n656), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G85), .A2(n650), .ZN(n651) );
  XNOR2_X1 U733 ( .A(KEYINPUT67), .B(n651), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n660), .A2(G60), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(G290) );
  NAND2_X1 U737 ( .A1(G49), .A2(n656), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n661), .A2(G87), .ZN(n662) );
  XOR2_X1 U742 ( .A(KEYINPUT79), .B(n662), .Z(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(G288) );
  XOR2_X1 U744 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n665) );
  XNOR2_X1 U745 ( .A(G305), .B(n665), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n666), .B(n676), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n715), .B(G166), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(n671) );
  XNOR2_X1 U749 ( .A(G290), .B(n994), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(G288), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n671), .B(n670), .ZN(n843) );
  XNOR2_X1 U752 ( .A(n843), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G868), .ZN(n674) );
  XOR2_X1 U754 ( .A(KEYINPUT83), .B(n674), .Z(n678) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U764 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G108), .A2(n684), .ZN(n842) );
  NAND2_X1 U766 ( .A1(G567), .A2(n842), .ZN(n685) );
  XNOR2_X1 U767 ( .A(n685), .B(KEYINPUT85), .ZN(n691) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n686) );
  XNOR2_X1 U769 ( .A(KEYINPUT22), .B(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n687), .A2(G96), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n688), .A2(G218), .ZN(n689) );
  XOR2_X1 U772 ( .A(n689), .B(KEYINPUT84), .Z(n841) );
  AND2_X1 U773 ( .A1(n841), .A2(G2106), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n691), .A2(n690), .ZN(G319) );
  INV_X1 U775 ( .A(G319), .ZN(n910) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U777 ( .A1(n910), .A2(n692), .ZN(n840) );
  NAND2_X1 U778 ( .A1(G36), .A2(n840), .ZN(n693) );
  XNOR2_X1 U779 ( .A(n693), .B(KEYINPUT86), .ZN(G176) );
  AND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n793) );
  NAND2_X1 U781 ( .A1(n795), .A2(n793), .ZN(n728) );
  INV_X1 U782 ( .A(n728), .ZN(n722) );
  INV_X1 U783 ( .A(n722), .ZN(n739) );
  NAND2_X1 U784 ( .A1(n739), .A2(G1341), .ZN(n697) );
  INV_X1 U785 ( .A(G1996), .ZN(n949) );
  NOR2_X1 U786 ( .A1(n728), .A2(n949), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n698), .A2(n994), .ZN(n699) );
  XOR2_X1 U790 ( .A(n699), .B(KEYINPUT64), .Z(n706) );
  OR2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n704) );
  AND2_X1 U792 ( .A1(n722), .A2(G2067), .ZN(n700) );
  XOR2_X1 U793 ( .A(n700), .B(KEYINPUT96), .Z(n702) );
  NAND2_X1 U794 ( .A1(n739), .A2(G1348), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n722), .A2(G2072), .ZN(n709) );
  XNOR2_X1 U800 ( .A(n709), .B(KEYINPUT27), .ZN(n711) );
  INV_X1 U801 ( .A(G1956), .ZN(n968) );
  NOR2_X1 U802 ( .A1(n968), .A2(n722), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U807 ( .A(n716), .B(KEYINPUT28), .Z(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U809 ( .A1(n722), .A2(G1961), .ZN(n721) );
  XNOR2_X1 U810 ( .A(n721), .B(KEYINPUT95), .ZN(n724) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NAND2_X1 U812 ( .A1(n722), .A2(n956), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n733) );
  NAND2_X1 U814 ( .A1(G171), .A2(n733), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U816 ( .A1(G8), .A2(n728), .ZN(n778) );
  NOR2_X1 U817 ( .A1(n778), .A2(G1966), .ZN(n727) );
  XNOR2_X1 U818 ( .A(n727), .B(KEYINPUT94), .ZN(n748) );
  NOR2_X1 U819 ( .A1(n728), .A2(G2084), .ZN(n750) );
  XNOR2_X1 U820 ( .A(n750), .B(KEYINPUT93), .ZN(n729) );
  NAND2_X1 U821 ( .A1(G8), .A2(n729), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n748), .A2(n730), .ZN(n731) );
  XOR2_X1 U823 ( .A(KEYINPUT30), .B(n731), .Z(n732) );
  NOR2_X1 U824 ( .A1(G168), .A2(n732), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G171), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n747) );
  NAND2_X1 U829 ( .A1(n747), .A2(G286), .ZN(n744) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n778), .ZN(n741) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n745), .A2(G8), .ZN(n746) );
  INV_X1 U836 ( .A(n770), .ZN(n755) );
  XNOR2_X1 U837 ( .A(KEYINPUT97), .B(n747), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n753) );
  XOR2_X1 U839 ( .A(KEYINPUT93), .B(n750), .Z(n751) );
  NAND2_X1 U840 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n769) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NAND2_X1 U843 ( .A1(n769), .A2(n1000), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n762) );
  INV_X1 U845 ( .A(n1000), .ZN(n757) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n763), .A2(n756), .ZN(n1004) );
  OR2_X1 U849 ( .A1(n757), .A2(n1004), .ZN(n758) );
  OR2_X1 U850 ( .A1(n778), .A2(n758), .ZN(n760) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n1007) );
  NAND2_X1 U854 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n520), .A2(n765), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT98), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n767) );
  XOR2_X1 U858 ( .A(KEYINPUT99), .B(n767), .Z(n768) );
  NAND2_X1 U859 ( .A1(n768), .A2(G8), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n778), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n780) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U865 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n817) );
  NAND2_X1 U868 ( .A1(G128), .A2(n891), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G116), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT35), .ZN(n791) );
  XNOR2_X1 U872 ( .A(KEYINPUT89), .B(KEYINPUT34), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n895), .A2(G140), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT88), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G104), .A2(n894), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n789), .B(n788), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT36), .B(n792), .Z(n907) );
  XNOR2_X1 U880 ( .A(G2067), .B(KEYINPUT37), .ZN(n829) );
  OR2_X1 U881 ( .A1(n907), .A2(n829), .ZN(n924) );
  INV_X1 U882 ( .A(n793), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U884 ( .A(KEYINPUT87), .B(n796), .Z(n831) );
  INV_X1 U885 ( .A(n831), .ZN(n815) );
  NOR2_X1 U886 ( .A1(n924), .A2(n815), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n797), .B(KEYINPUT90), .ZN(n827) );
  NAND2_X1 U888 ( .A1(G95), .A2(n894), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G119), .A2(n891), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G131), .A2(n895), .ZN(n800) );
  XNOR2_X1 U892 ( .A(KEYINPUT91), .B(n800), .ZN(n801) );
  NOR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G107), .A2(n781), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n889) );
  AND2_X1 U896 ( .A1(n889), .A2(G1991), .ZN(n814) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n806) );
  NAND2_X1 U898 ( .A1(G105), .A2(n894), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n806), .B(n805), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G141), .A2(n895), .ZN(n808) );
  NAND2_X1 U901 ( .A1(G129), .A2(n891), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G117), .A2(n781), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n888) );
  AND2_X1 U906 ( .A1(n888), .A2(G1996), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n921) );
  NOR2_X1 U908 ( .A1(n921), .A2(n815), .ZN(n823) );
  OR2_X1 U909 ( .A1(n827), .A2(n823), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT100), .ZN(n820) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n1006) );
  NAND2_X1 U913 ( .A1(n1006), .A2(n831), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n834) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n888), .ZN(n918) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n889), .ZN(n923) );
  NOR2_X1 U918 ( .A1(n821), .A2(n923), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n918), .A2(n824), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT39), .B(n825), .Z(n826) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n828), .B(KEYINPUT101), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n907), .A2(n829), .ZN(n938) );
  NAND2_X1 U925 ( .A1(n830), .A2(n938), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XOR2_X1 U941 ( .A(KEYINPUT112), .B(n843), .Z(n845) );
  XNOR2_X1 U942 ( .A(G171), .B(G286), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n993), .B(n846), .ZN(n847) );
  NOR2_X1 U945 ( .A1(G37), .A2(n847), .ZN(G397) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2100), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G2096), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1981), .B(G1956), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1961), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n867) );
  XOR2_X1 U958 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1991), .B(KEYINPUT106), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(G1976), .B(G1971), .Z(n861) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1986), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT107), .B(G2474), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(G229) );
  XOR2_X1 U968 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n869) );
  NAND2_X1 U969 ( .A1(G124), .A2(n891), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n870), .B(KEYINPUT108), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n894), .A2(G100), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G136), .A2(n895), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G112), .A2(n781), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U977 ( .A1(n876), .A2(n875), .ZN(G162) );
  XOR2_X1 U978 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n886) );
  NAND2_X1 U979 ( .A1(G103), .A2(n894), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G139), .A2(n895), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G127), .A2(n891), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G115), .A2(n781), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  XNOR2_X1 U986 ( .A(KEYINPUT110), .B(n882), .ZN(n883) );
  NOR2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n931) );
  XNOR2_X1 U988 ( .A(n931), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(n888), .B(n887), .Z(n906) );
  XNOR2_X1 U991 ( .A(G162), .B(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n890), .B(n920), .ZN(n902) );
  NAND2_X1 U993 ( .A1(G130), .A2(n891), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G118), .A2(n781), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G106), .A2(n894), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G142), .A2(n895), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(KEYINPUT45), .B(n898), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G164), .B(G160), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n910), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n915), .A2(G395), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1016 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1029) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n1020) );
  XOR2_X1 U1018 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n941) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n919), .Z(n930) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(n928), .B(KEYINPUT114), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G164), .B(G2078), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT115), .B(n935), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n941), .B(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n1020), .A2(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1039 ( .A(KEYINPUT117), .B(G2090), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(G35), .ZN(n965) );
  XOR2_X1 U1041 ( .A(G34), .B(KEYINPUT121), .Z(n946) );
  XNOR2_X1 U1042 ( .A(G2084), .B(KEYINPUT54), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n946), .B(n945), .ZN(n963) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G32), .B(n949), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n950), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(G25), .B(G1991), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n951), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G27), .B(n956), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(KEYINPUT119), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n960), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n1021) );
  NOR2_X1 U1060 ( .A1(G29), .A2(KEYINPUT55), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n1021), .A2(n966), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n967), .ZN(n1025) );
  XOR2_X1 U1063 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n990) );
  XNOR2_X1 U1064 ( .A(G20), .B(n968), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n973) );
  XNOR2_X1 U1070 ( .A(G4), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G5), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n988) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(G1976), .B(G23), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1078 ( .A(KEYINPUT124), .B(n981), .Z(n983) );
  XNOR2_X1 U1079 ( .A(G1986), .B(G24), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1081 ( .A(KEYINPUT58), .B(n984), .Z(n986) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G21), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n990), .B(n989), .ZN(n992) );
  XOR2_X1 U1086 ( .A(KEYINPUT123), .B(G16), .Z(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n1018) );
  XOR2_X1 U1088 ( .A(G16), .B(KEYINPUT56), .Z(n1015) );
  XNOR2_X1 U1089 ( .A(G1348), .B(n993), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G301), .B(G1961), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n994), .B(G1341), .ZN(n995) );
  NOR2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n1013) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(G1956), .B(G299), .ZN(n1001) );
  NOR2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1102 ( .A(n1009), .B(KEYINPUT57), .ZN(n1010) );
  NAND2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(KEYINPUT122), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1019), .ZN(n1023) );
  OR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(n1029), .B(n1028), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

