//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  XOR2_X1   g000(.A(KEYINPUT87), .B(G104), .Z(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G237), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT73), .ZN(new_n195));
  OAI211_X1 g009(.A(G214), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(KEYINPUT73), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(G237), .ZN(new_n200));
  AOI21_X1  g014(.A(G953), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(G143), .A3(G214), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT18), .A2(G131), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n203), .B(KEYINPUT86), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT65), .A2(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT65), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(new_n210), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n198), .A2(new_n202), .ZN(new_n218));
  INV_X1    g032(.A(new_n203), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT85), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT19), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n210), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n215), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT65), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n227), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n196), .A2(new_n197), .ZN(new_n235));
  AOI21_X1  g049(.A(G143), .B1(new_n201), .B2(G214), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT67), .A2(G131), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT67), .A2(G131), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n235), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n237), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n198), .A2(new_n240), .A3(new_n202), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n234), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n190), .B1(new_n224), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n205), .A2(new_n216), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n222), .B1(new_n218), .B2(new_n219), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT85), .B(new_n203), .C1(new_n198), .C2(new_n202), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n248), .A3(new_n241), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n225), .A2(new_n226), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n227), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n240), .B1(new_n198), .B2(new_n202), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n247), .A2(new_n255), .A3(new_n189), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n243), .A2(new_n256), .ZN(new_n257));
  NOR3_X1   g071(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n247), .A2(new_n255), .A3(new_n189), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n239), .A2(new_n241), .ZN(new_n262));
  INV_X1    g076(.A(new_n227), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n210), .B(KEYINPUT19), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n213), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n189), .B1(new_n247), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n260), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G475), .A2(G902), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n243), .A2(KEYINPUT88), .A3(new_n256), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n259), .B1(new_n271), .B2(KEYINPUT20), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n191), .A2(G952), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(G234), .B2(G237), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n275), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT21), .B(G898), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G122), .ZN(new_n279));
  OR3_X1    g093(.A1(new_n279), .A2(KEYINPUT14), .A3(G116), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G122), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(G116), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n283), .A3(KEYINPUT90), .A4(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(G107), .C1(KEYINPUT90), .C2(new_n280), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n284), .A2(new_n282), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G128), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n290), .A2(KEYINPUT89), .A3(G143), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT89), .B1(new_n290), .B2(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n290), .A2(G143), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G134), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n293), .A2(G134), .A3(new_n294), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n286), .B(new_n289), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  INV_X1    g114(.A(G217), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(G953), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT91), .ZN(new_n303));
  INV_X1    g117(.A(new_n298), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n294), .B(KEYINPUT13), .ZN(new_n305));
  OAI21_X1  g119(.A(G134), .B1(new_n305), .B2(new_n293), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n287), .B(new_n288), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n299), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n303), .B1(new_n299), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n275), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G478), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(KEYINPUT15), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G475), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n189), .B1(new_n247), .B2(new_n255), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n261), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n275), .ZN(new_n318));
  NOR4_X1   g132(.A1(new_n272), .A2(new_n278), .A3(new_n314), .A4(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n296), .B2(G137), .ZN(new_n323));
  INV_X1    g137(.A(G137), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT11), .A3(G134), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n324), .A2(G134), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n327), .A2(new_n238), .A3(new_n237), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n325), .ZN(new_n331));
  OR2_X1    g145(.A1(KEYINPUT67), .A2(G131), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n296), .A2(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT67), .A2(G131), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT68), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n326), .A2(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n197), .A2(G146), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT1), .ZN(new_n342));
  OAI21_X1  g156(.A(G128), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n211), .A2(new_n212), .A3(new_n197), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT66), .B1(new_n215), .B2(G143), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n197), .A3(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n343), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n231), .A2(G143), .A3(new_n232), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n290), .A2(KEYINPUT1), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n347), .A3(new_n345), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n288), .A2(G104), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G107), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n359), .A2(KEYINPUT3), .B1(new_n288), .B2(G104), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n361));
  OAI22_X1  g175(.A1(KEYINPUT79), .A2(new_n361), .B1(new_n356), .B2(G107), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n288), .A3(KEYINPUT3), .A4(G104), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n358), .B1(new_n364), .B2(new_n354), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n290), .B1(new_n350), .B2(KEYINPUT1), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n341), .B1(new_n233), .B2(new_n197), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n352), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n365), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n340), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT12), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT72), .B(new_n352), .C1(new_n367), .C2(new_n368), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n376), .B(new_n358), .C1(new_n364), .C2(new_n354), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n353), .A2(new_n365), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n376), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n344), .A2(new_n348), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n341), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n213), .B2(G143), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT0), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n290), .A3(KEYINPUT64), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(KEYINPUT0), .B2(G128), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n381), .A2(new_n383), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n362), .A2(new_n363), .ZN(new_n392));
  INV_X1    g206(.A(new_n360), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G101), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT4), .B1(new_n394), .B2(G101), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n364), .A2(new_n354), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n391), .B(new_n396), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n330), .A2(new_n336), .B1(new_n338), .B2(G131), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n378), .A2(new_n380), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n191), .A2(G227), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(new_n340), .C1(new_n366), .C2(new_n370), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n372), .A2(new_n401), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n378), .A2(new_n380), .A3(new_n399), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n340), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n410), .B2(new_n401), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n408), .B1(new_n411), .B2(KEYINPUT81), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n372), .A2(new_n401), .A3(new_n407), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT80), .B(G469), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n275), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n404), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT10), .B1(new_n353), .B2(new_n365), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT4), .B(new_n354), .C1(new_n392), .C2(new_n393), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n394), .A2(G101), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n395), .B1(new_n364), .B2(new_n354), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n425), .B2(new_n391), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n400), .B1(new_n426), .B2(new_n378), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n400), .A2(new_n378), .A3(new_n380), .A4(new_n399), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n405), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G469), .B1(new_n430), .B2(G902), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n321), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n281), .B2(G119), .ZN(new_n436));
  INV_X1    g250(.A(G119), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT71), .A3(G116), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n281), .A2(G119), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT2), .B(G113), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n396), .C1(new_n397), .C2(new_n398), .ZN(new_n443));
  INV_X1    g257(.A(G113), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n445));
  NOR2_X1   g259(.A1(new_n281), .A2(G119), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n440), .B2(new_n445), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n440), .A2(new_n441), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n365), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n450), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n381), .A2(new_n383), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n385), .A2(new_n390), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G125), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n208), .B(new_n352), .C1(new_n367), .C2(new_n368), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n391), .A2(new_n208), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n463), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n470), .A2(new_n473), .A3(new_n462), .ZN(new_n476));
  OAI22_X1  g290(.A1(new_n458), .A2(new_n460), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n447), .B1(new_n478), .B2(new_n440), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n449), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n365), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n451), .B(KEYINPUT8), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n448), .A2(new_n449), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n481), .B(new_n482), .C1(new_n365), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n485));
  INV_X1    g299(.A(new_n469), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n472), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n452), .A3(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n470), .A2(new_n473), .A3(new_n485), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n275), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n477), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n492), .ZN(new_n494));
  INV_X1    g308(.A(new_n476), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n462), .B1(new_n470), .B2(new_n473), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n495), .A2(new_n496), .B1(new_n457), .B2(new_n459), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n497), .B2(new_n490), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n434), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n319), .A2(new_n432), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n296), .A2(KEYINPUT69), .A3(G137), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT69), .B1(new_n296), .B2(G137), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n333), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G131), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n369), .A2(new_n337), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n506), .A2(KEYINPUT70), .B1(new_n340), .B2(new_n391), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n330), .A2(new_n336), .B1(G131), .B2(new_n504), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n369), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT30), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n374), .A2(new_n508), .A3(new_n375), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT30), .B1(new_n400), .B2(new_n467), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n442), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n374), .A2(new_n508), .A3(new_n375), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n340), .A2(new_n391), .ZN(new_n517));
  INV_X1    g331(.A(new_n442), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n201), .A2(G210), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT27), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT74), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n527), .C1(new_n511), .C2(new_n514), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n516), .A2(new_n532), .A3(new_n517), .A4(new_n518), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n506), .A2(KEYINPUT70), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n510), .A3(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n442), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n513), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n518), .B1(new_n541), .B2(new_n516), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n524), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n530), .A2(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n529), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G472), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n519), .B1(new_n511), .B2(new_n514), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n530), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n534), .A2(new_n523), .A3(new_n537), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n518), .B1(new_n516), .B2(new_n517), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n531), .B2(new_n533), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n530), .A2(new_n555), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n552), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n547), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n529), .B2(new_n545), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(KEYINPUT32), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT75), .B1(new_n564), .B2(KEYINPUT32), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n551), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n290), .A2(KEYINPUT23), .A3(G119), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n437), .A2(G128), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n437), .A2(G128), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(KEYINPUT23), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  XNOR2_X1  g386(.A(G119), .B(G128), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n571), .A2(G110), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(G146), .B1(new_n225), .B2(new_n226), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n263), .B2(new_n575), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n571), .A2(G110), .B1(new_n572), .B2(new_n573), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n227), .A3(new_n214), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n578), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT77), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n301), .B1(G234), .B2(new_n275), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n275), .A3(new_n585), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n584), .A2(KEYINPUT25), .A3(new_n275), .A4(new_n585), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(KEYINPUT76), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n597), .A3(new_n593), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n588), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n501), .A2(new_n567), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n546), .A2(new_n275), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(new_n432), .A3(new_n548), .A4(new_n601), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n318), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n271), .A2(KEYINPUT20), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n259), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n310), .A2(KEYINPUT93), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n309), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n310), .A2(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n309), .B2(new_n310), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT92), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(KEYINPUT92), .B(new_n612), .C1(new_n309), .C2(new_n310), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n312), .A2(G902), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n615), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n311), .A2(new_n312), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n610), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n278), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n499), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n607), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n271), .A2(KEYINPUT20), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT20), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n268), .A2(new_n632), .A3(new_n270), .A4(new_n269), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n608), .A3(new_n314), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n607), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT94), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n583), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n579), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n589), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n599), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n599), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n599), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n599), .A2(new_n642), .A3(new_n645), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(KEYINPUT96), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n605), .A3(new_n548), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(new_n500), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n276), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n274), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n634), .A2(new_n608), .A3(new_n314), .A4(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n652), .B2(new_n648), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n432), .A2(new_n499), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n567), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n493), .A2(new_n498), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT38), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n610), .A2(new_n314), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n650), .A2(new_n651), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n669), .A2(new_n670), .A3(new_n434), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n558), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n519), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n530), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n525), .A2(new_n528), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n275), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n564), .A2(KEYINPUT32), .B1(new_n677), .B2(G472), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n551), .A2(new_n678), .A3(new_n566), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n662), .B(KEYINPUT39), .Z(new_n680));
  AOI211_X1 g494(.A(new_n321), .B(new_n680), .C1(new_n419), .C2(new_n431), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT40), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  OAI211_X1 g498(.A(new_n623), .B(new_n662), .C1(new_n272), .C2(new_n318), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n652), .B2(new_n648), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n567), .A2(new_n665), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT98), .B(G146), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G48));
  AND2_X1   g503(.A1(new_n567), .A2(new_n601), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n404), .B1(new_n427), .B2(new_n428), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n691), .A2(new_n414), .B1(new_n413), .B2(new_n405), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n408), .A2(KEYINPUT81), .ZN(new_n693));
  OAI211_X1 g507(.A(KEYINPUT99), .B(new_n275), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n412), .B2(new_n415), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n419), .B(new_n320), .C1(new_n695), .C2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n624), .A3(new_n626), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n690), .A2(KEYINPUT100), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n698), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n567), .A3(new_n627), .A4(new_n601), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n701), .A2(new_n567), .A3(new_n636), .A4(new_n601), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND2_X1  g523(.A1(new_n567), .A2(new_n653), .ZN(new_n710));
  AOI211_X1 g524(.A(G902), .B(new_n417), .C1(new_n412), .C2(new_n415), .ZN(new_n711));
  INV_X1    g525(.A(new_n697), .ZN(new_n712));
  INV_X1    g526(.A(G469), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n696), .B2(KEYINPUT99), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n320), .A3(new_n499), .A4(new_n319), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n437), .ZN(G21));
  NOR3_X1   g532(.A1(new_n698), .A2(new_n626), .A3(new_n670), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n552), .B1(new_n546), .B2(new_n275), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n559), .A2(new_n523), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n529), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT101), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n543), .A2(new_n544), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n529), .A2(new_n725), .A3(new_n721), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n720), .B1(new_n727), .B2(new_n547), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n601), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n728), .B2(new_n601), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n719), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  INV_X1    g548(.A(new_n499), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n698), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n685), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n671), .A3(new_n728), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n548), .A2(new_n550), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n565), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n601), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n493), .A2(new_n498), .A3(new_n433), .ZN(new_n743));
  INV_X1    g557(.A(new_n320), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n419), .B2(new_n431), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n737), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT42), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n745), .A2(new_n743), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n567), .A2(new_n748), .A3(new_n601), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(G131), .Z(G33));
  INV_X1    g566(.A(new_n663), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n567), .A2(new_n748), .A3(new_n753), .A4(new_n601), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NOR2_X1   g569(.A1(new_n272), .A2(new_n318), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n623), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n671), .C1(new_n564), .C2(new_n720), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n743), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n430), .A2(KEYINPUT45), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n420), .A2(new_n769), .A3(new_n429), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n419), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n320), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n680), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n765), .A2(new_n767), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT104), .B(G137), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  NOR4_X1   g596(.A1(new_n567), .A2(new_n601), .A3(new_n685), .A4(new_n766), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT106), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(KEYINPUT106), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n711), .B1(new_n773), .B2(new_n774), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n744), .B(new_n787), .C1(new_n788), .C2(new_n776), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n777), .B2(new_n320), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n784), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n206), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n794));
  NOR2_X1   g608(.A1(G952), .A2(G953), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT116), .Z(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n698), .A2(new_n661), .A3(new_n766), .ZN(new_n798));
  INV_X1    g612(.A(new_n679), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n610), .A2(new_n623), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n601), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n727), .A2(new_n547), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n605), .A3(new_n671), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n798), .A2(new_n762), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n715), .A2(new_n321), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n766), .B1(new_n791), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n762), .A2(new_n274), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n601), .A3(new_n605), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT102), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n810), .B2(new_n730), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n698), .A2(KEYINPUT111), .A3(new_n433), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT111), .B1(new_n698), .B2(new_n433), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n814), .A2(new_n669), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n817), .B2(KEYINPUT112), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n819), .B(KEYINPUT50), .C1(new_n811), .C2(new_n816), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n812), .B(KEYINPUT51), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  INV_X1    g636(.A(new_n808), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n731), .B2(new_n732), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n669), .A3(new_n815), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT50), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n813), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT51), .A4(new_n812), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n804), .A2(new_n742), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n798), .A2(new_n601), .A3(new_n799), .ZN(new_n836));
  INV_X1    g650(.A(new_n624), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n273), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT114), .B1(new_n811), .B2(new_n736), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n811), .A2(KEYINPUT114), .A3(new_n736), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n835), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n812), .B1(new_n818), .B2(new_n820), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n832), .A2(new_n833), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n833), .B1(new_n832), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n610), .A2(new_n499), .A3(new_n314), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n662), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n649), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n679), .A2(new_n745), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n567), .B(new_n665), .C1(new_n664), .C2(new_n686), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n738), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n708), .B1(new_n710), .B2(new_n716), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n705), .A2(new_n858), .A3(new_n733), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT107), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n501), .A2(new_n567), .A3(new_n601), .ZN(new_n861));
  INV_X1    g675(.A(new_n623), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n610), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n314), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n756), .A2(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n434), .B(new_n278), .C1(new_n493), .C2(new_n498), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n606), .A2(new_n867), .B1(new_n654), .B2(new_n500), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n860), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n867), .A2(new_n606), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n655), .A3(new_n602), .A4(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n314), .A2(new_n850), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n608), .A2(new_n743), .A3(new_n634), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n567), .A2(new_n874), .A3(new_n432), .A4(new_n653), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n754), .B(new_n875), .C1(new_n803), .C2(new_n746), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n751), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n856), .A2(new_n859), .A3(new_n872), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n857), .B1(new_n704), .B2(new_n700), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n872), .A3(new_n877), .A4(new_n733), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n852), .A2(new_n687), .A3(KEYINPUT52), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n715), .A2(new_n320), .A3(new_n499), .A4(new_n737), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n666), .B(KEYINPUT108), .C1(new_n803), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT108), .B1(new_n738), .B2(new_n666), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n853), .A2(new_n852), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n803), .A2(new_n885), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n855), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT109), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT109), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n854), .A2(new_n894), .A3(new_n855), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT110), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT110), .A4(new_n895), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n883), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n881), .B1(new_n900), .B2(KEYINPUT53), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n872), .A4(new_n877), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n854), .A2(new_n894), .A3(new_n855), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n894), .B1(new_n854), .B2(new_n855), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT110), .B1(new_n906), .B2(new_n889), .ZN(new_n907));
  INV_X1    g721(.A(new_n899), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT54), .B1(new_n878), .B2(new_n879), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n901), .A2(KEYINPUT54), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n797), .B1(new_n847), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n715), .B(KEYINPUT49), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n610), .A2(new_n862), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n600), .A2(new_n321), .A3(new_n434), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n799), .A2(new_n669), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n794), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n917), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n909), .A2(new_n910), .ZN(new_n920));
  INV_X1    g734(.A(new_n883), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n907), .B2(new_n908), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n880), .B1(new_n922), .B2(new_n879), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n925), .A2(new_n846), .A3(new_n845), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT117), .B(new_n919), .C1(new_n926), .C2(new_n797), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n918), .A2(new_n927), .ZN(G75));
  AOI21_X1  g742(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n854), .B(KEYINPUT52), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n879), .B1(new_n883), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n275), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n458), .A2(new_n460), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n495), .A3(new_n496), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n477), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  AND3_X1   g754(.A1(new_n935), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n935), .B2(new_n936), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n191), .A2(G952), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G51));
  NAND3_X1  g758(.A1(new_n909), .A2(KEYINPUT118), .A3(new_n910), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n931), .A2(new_n924), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n929), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT54), .B1(new_n929), .B2(new_n932), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n772), .B(KEYINPUT57), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n416), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n933), .A2(new_n275), .A3(new_n771), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(G54));
  INV_X1    g769(.A(new_n943), .ZN(new_n956));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n934), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n268), .A2(new_n270), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT119), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  AND4_X1   g776(.A1(KEYINPUT119), .A2(new_n934), .A3(new_n960), .A4(new_n957), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G60));
  NAND3_X1  g778(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT59), .Z(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT120), .B1(new_n950), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n950), .A2(KEYINPUT120), .A3(new_n968), .ZN(new_n970));
  INV_X1    g784(.A(new_n965), .ZN(new_n971));
  INV_X1    g785(.A(new_n967), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n925), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n974));
  OAI22_X1  g788(.A1(new_n969), .A2(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n965), .B1(new_n911), .B2(new_n967), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n956), .B1(new_n976), .B2(KEYINPUT121), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G63));
  INV_X1    g792(.A(new_n933), .ZN(new_n979));
  XNOR2_X1  g793(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n301), .A2(new_n275), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n587), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n979), .A2(new_n644), .A3(new_n982), .ZN(new_n985));
  NOR2_X1   g799(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n943), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G66));
  INV_X1    g804(.A(new_n277), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n191), .B1(new_n991), .B2(G224), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n859), .A2(new_n872), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n191), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n937), .B1(G898), .B2(new_n191), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n994), .B(new_n995), .Z(G69));
  OAI21_X1  g810(.A(new_n540), .B1(new_n512), .B2(new_n513), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n229), .B(KEYINPUT124), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n887), .A2(new_n888), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n687), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n683), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n780), .A2(new_n792), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n863), .A2(new_n865), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n690), .A2(new_n681), .A3(new_n743), .A4(new_n1006), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1003), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n999), .B1(new_n1009), .B2(new_n191), .ZN(new_n1010));
  INV_X1    g824(.A(new_n779), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n849), .A2(new_n741), .A3(new_n601), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n754), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n1012), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1014), .A2(new_n751), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1017), .A2(G953), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G900), .A2(G953), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n1018), .A2(new_n999), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(G72));
  INV_X1    g837(.A(new_n553), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1024), .A2(new_n530), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n993), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1003), .A2(new_n1027), .A3(new_n1004), .A4(new_n1008), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  AOI21_X1  g844(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT126), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n525), .A2(new_n554), .A3(new_n528), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n901), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1030), .B1(new_n1017), .B2(new_n993), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT127), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1024), .A2(new_n530), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n956), .B(new_n1034), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1032), .A2(new_n1038), .ZN(G57));
endmodule


