//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(KEYINPUT87), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(KEYINPUT87), .B2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT14), .B(G29gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G1gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G1gat), .B2(new_n217), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G8gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n214), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n223), .A2(KEYINPUT18), .A3(new_n224), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n214), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n224), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n229), .A2(new_n242), .A3(new_n230), .A4(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G127gat), .A2(G134gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(G127gat), .A2(G134gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(G113gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G120gat), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n248), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n258));
  INV_X1    g057(.A(G155gat), .ZN(new_n259));
  INV_X1    g058(.A(G162gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G148gat), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n261), .A2(new_n262), .B1(new_n264), .B2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g064(.A(G148gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G141gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(G148gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(G141gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n258), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n265), .A2(new_n270), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n254), .B2(G120gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n252), .A3(G113gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n280), .A3(new_n255), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n246), .B2(new_n247), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n277), .A2(new_n281), .A3(new_n249), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n257), .A2(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n262), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n270), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G141gat), .B(G148gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n275), .B1(new_n292), .B2(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n257), .A2(new_n276), .A3(KEYINPUT4), .A4(new_n284), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n287), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT5), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n287), .A2(new_n298), .A3(new_n301), .A4(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n294), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n305), .B2(new_n285), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT0), .ZN(new_n309));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n302), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(new_n307), .ZN(new_n316));
  INV_X1    g115(.A(new_n311), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(G211gat), .A2(G218gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(G197gat), .A2(G204gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G197gat), .A2(G204gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n320), .A2(KEYINPUT22), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G197gat), .B(G204gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  INV_X1    g129(.A(G211gat), .ZN(new_n331));
  INV_X1    g130(.A(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT26), .ZN(new_n338));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n339), .C1(new_n342), .C2(new_n337), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n348), .B2(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT28), .A4(new_n352), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n343), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n358), .A2(new_n340), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n364), .A2(new_n365), .B1(new_n339), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n367), .B2(KEYINPUT65), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n339), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n369), .A2(KEYINPUT65), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n357), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n362), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n356), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(KEYINPUT29), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n377), .B(new_n356), .C1(new_n372), .C2(new_n374), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n336), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n372), .A2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(new_n356), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n376), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n384), .B(new_n335), .C1(new_n375), .C2(new_n378), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n379), .A2(new_n380), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n335), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n398), .A3(new_n393), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n319), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n297), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n297), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n336), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n327), .B2(new_n334), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n294), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n294), .B2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(new_n336), .ZN(new_n412));
  INV_X1    g211(.A(new_n296), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n294), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT79), .B1(new_n415), .B2(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  INV_X1    g216(.A(new_n409), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n417), .B(new_n418), .C1(new_n412), .C2(new_n414), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n411), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n411), .C1(new_n416), .C2(new_n419), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT82), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n422), .A3(new_n427), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT78), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT31), .B(G50gat), .Z(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n426), .A2(new_n431), .A3(new_n435), .A4(new_n428), .ZN(new_n438));
  XNOR2_X1  g237(.A(G15gat), .B(G43gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n382), .A2(new_n383), .ZN(new_n442));
  INV_X1    g241(.A(new_n288), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G227gat), .ZN(new_n445));
  INV_X1    g244(.A(G233gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n375), .A2(new_n288), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n441), .B1(new_n449), .B2(KEYINPUT32), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n444), .A2(new_n448), .ZN(new_n454));
  INV_X1    g253(.A(new_n447), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT72), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n447), .B1(new_n444), .B2(new_n448), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n441), .A2(KEYINPUT71), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n441), .A2(KEYINPUT71), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT33), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT32), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n453), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n453), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n400), .A2(new_n437), .A3(new_n438), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n472), .A3(KEYINPUT35), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n437), .A2(new_n468), .A3(new_n438), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  INV_X1    g275(.A(new_n397), .ZN(new_n477));
  INV_X1    g276(.A(new_n399), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n397), .A2(KEYINPUT83), .A3(new_n399), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n319), .A2(KEYINPUT35), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n471), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n300), .A2(new_n301), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n305), .A2(new_n301), .A3(new_n285), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(KEYINPUT39), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n317), .C1(KEYINPUT39), .C2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n312), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n479), .A2(new_n493), .A3(new_n480), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n319), .A2(new_n394), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n395), .A2(KEYINPUT37), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n396), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n390), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT38), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n381), .B2(new_n385), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n501), .B2(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n497), .A2(new_n502), .A3(new_n506), .A4(new_n503), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n495), .A2(new_n500), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n437), .A2(new_n438), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n468), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n468), .B1(new_n515), .B2(new_n513), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n400), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n511), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n245), .B1(new_n484), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G127gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n222), .B1(new_n527), .B2(new_n526), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(new_n259), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT90), .ZN(new_n543));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT8), .ZN(new_n552));
  AND2_X1   g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT91), .B(G85gat), .Z(new_n554));
  OAI221_X1 g353(.A(new_n551), .B1(new_n552), .B2(new_n553), .C1(G92gat), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT92), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n555), .A2(new_n557), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n216), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n558), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(new_n225), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n549), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n547), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n563), .A2(new_n566), .A3(new_n549), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n570), .A2(new_n568), .A3(new_n571), .A4(new_n547), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n541), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n558), .A3(new_n526), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n580));
  INV_X1    g379(.A(new_n526), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n561), .A3(new_n559), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n565), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n582), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n578), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n521), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n319), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(G1gat), .Z(G1324gat));
  INV_X1    g399(.A(new_n481), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n521), .A2(new_n601), .A3(new_n596), .ZN(new_n602));
  AND2_X1   g401(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT42), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n602), .A2(G8gat), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n608), .B(new_n609), .C1(new_n606), .C2(new_n605), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n597), .B2(new_n517), .ZN(new_n611));
  INV_X1    g410(.A(new_n468), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(G15gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n597), .B2(new_n613), .ZN(G1326gat));
  NOR2_X1   g413(.A1(new_n597), .A2(new_n510), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT43), .B(G22gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(G1327gat));
  AOI21_X1  g416(.A(new_n575), .B1(new_n484), .B2(new_n520), .ZN(new_n618));
  NAND2_X1  g417(.A1(KEYINPUT97), .A2(KEYINPUT44), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(KEYINPUT97), .A2(KEYINPUT44), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n541), .B(KEYINPUT96), .Z(new_n626));
  NOR4_X1   g425(.A1(new_n625), .A2(new_n245), .A3(new_n595), .A4(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(G29gat), .B1(new_n628), .B2(new_n598), .ZN(new_n629));
  INV_X1    g428(.A(new_n575), .ZN(new_n630));
  INV_X1    g429(.A(new_n541), .ZN(new_n631));
  INV_X1    g430(.A(new_n595), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n521), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n633), .A2(G29gat), .A3(new_n598), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT45), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(G1328gat));
  OAI21_X1  g435(.A(G36gat), .B1(new_n628), .B2(new_n481), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n633), .A2(G36gat), .A3(new_n481), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT46), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(G1329gat));
  NOR3_X1   g439(.A1(new_n633), .A2(G43gat), .A3(new_n612), .ZN(new_n641));
  INV_X1    g440(.A(new_n517), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n643), .B2(G43gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g444(.A1(new_n633), .A2(G50gat), .A3(new_n510), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n509), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(G50gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g448(.A1(new_n484), .A2(new_n520), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n576), .A2(new_n244), .A3(new_n632), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n598), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g453(.A(new_n652), .B(KEYINPUT98), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n481), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT99), .Z(new_n658));
  NOR2_X1   g457(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1333gat));
  NAND3_X1  g459(.A1(new_n655), .A2(G71gat), .A3(new_n642), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n652), .A2(new_n612), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n661), .B(KEYINPUT100), .C1(G71gat), .C2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(KEYINPUT100), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g464(.A1(new_n655), .A2(new_n509), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT101), .B(G78gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1335gat));
  NOR2_X1   g467(.A1(new_n541), .A2(new_n244), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n630), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT51), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n618), .A2(KEYINPUT51), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR4_X1    g474(.A1(new_n598), .A2(new_n675), .A3(new_n554), .A4(new_n632), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n541), .A2(new_n244), .A3(new_n632), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n618), .A2(new_n623), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n575), .B(new_n621), .C1(new_n484), .C2(new_n520), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n624), .A2(new_n682), .A3(new_n677), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n683), .A3(new_n319), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n554), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n676), .A2(new_n685), .ZN(G1336gat));
  OAI211_X1 g485(.A(new_n601), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT104), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n624), .A2(new_n689), .A3(new_n601), .A4(new_n677), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n690), .A3(G92gat), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n632), .B1(new_n672), .B2(new_n673), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n481), .A2(G92gat), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT52), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(KEYINPUT105), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n694), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND4_X1   g497(.A1(KEYINPUT51), .A2(new_n650), .A3(new_n630), .A4(new_n669), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT51), .B1(new_n618), .B2(new_n669), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n595), .B(new_n693), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n674), .A2(KEYINPUT103), .A3(new_n595), .A4(new_n693), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n681), .A2(new_n683), .A3(new_n601), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(G92gat), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n695), .B(new_n698), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n706), .A2(G92gat), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT52), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n695), .A4(new_n698), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(G1337gat));
  NAND3_X1  g514(.A1(new_n681), .A2(new_n683), .A3(new_n642), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G99gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n632), .A2(new_n612), .A3(G99gat), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT108), .Z(new_n722));
  OAI22_X1  g521(.A1(new_n719), .A2(new_n720), .B1(new_n675), .B2(new_n722), .ZN(G1338gat));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n681), .A2(new_n683), .A3(new_n509), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G106gat), .ZN(new_n726));
  INV_X1    g525(.A(G106gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n692), .A2(new_n727), .A3(new_n509), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n732));
  OAI21_X1  g531(.A(G106gat), .B1(new_n680), .B2(new_n510), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT111), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n730), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n735), .A3(new_n736), .ZN(G1339gat));
  NAND2_X1  g536(.A1(new_n596), .A2(new_n245), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n583), .A2(new_n578), .A3(new_n584), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n592), .A2(KEYINPUT54), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n590), .B1(new_n585), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(KEYINPUT55), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n594), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n244), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n232), .A2(new_n233), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n239), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n243), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n595), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n575), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n574), .A3(new_n573), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n749), .A2(new_n594), .A3(new_n744), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT112), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n745), .B1(new_n748), .B2(new_n747), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n630), .A4(new_n754), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n626), .B1(new_n764), .B2(KEYINPUT113), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n757), .A2(new_n766), .A3(new_n760), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n739), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n768), .A2(new_n598), .A3(new_n601), .A4(new_n474), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT115), .Z(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n254), .A3(new_n244), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n760), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n630), .B1(new_n750), .B2(new_n755), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT113), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n541), .B(KEYINPUT96), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n738), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n510), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT114), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n601), .A2(new_n598), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n468), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G113gat), .B1(new_n781), .B2(new_n245), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n782), .ZN(G1340gat));
  NAND3_X1  g582(.A1(new_n770), .A2(new_n252), .A3(new_n595), .ZN(new_n784));
  OAI21_X1  g583(.A(G120gat), .B1(new_n781), .B2(new_n632), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1341gat));
  OAI21_X1  g585(.A(G127gat), .B1(new_n781), .B2(new_n775), .ZN(new_n787));
  INV_X1    g586(.A(G127gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n788), .A3(new_n541), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1342gat));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  AOI21_X1  g590(.A(G134gat), .B1(new_n791), .B2(KEYINPUT56), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n769), .A2(new_n630), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(KEYINPUT56), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G134gat), .B1(new_n781), .B2(new_n575), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1343gat));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n777), .A2(new_n798), .A3(new_n509), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n517), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n747), .A2(new_n803), .A3(new_n748), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n747), .B2(new_n748), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT118), .B(new_n746), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n244), .ZN(new_n808));
  INV_X1    g607(.A(new_n806), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n804), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT118), .B1(new_n810), .B2(new_n746), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n755), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n772), .B1(new_n812), .B2(new_n575), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n738), .B1(new_n813), .B2(new_n541), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n798), .B1(new_n814), .B2(new_n509), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n802), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G141gat), .B1(new_n817), .B2(new_n245), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n768), .A2(new_n598), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n642), .A2(new_n510), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(KEYINPUT119), .A3(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n481), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n244), .A2(new_n263), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n818), .B(new_n819), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n822), .A2(new_n601), .A3(new_n827), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n818), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n830), .B2(new_n819), .ZN(G1344gat));
  OR2_X1    g630(.A1(new_n266), .A2(KEYINPUT59), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n816), .B2(new_n595), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n510), .A2(KEYINPUT57), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n812), .A2(new_n575), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n758), .A2(new_n759), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n541), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n837), .B2(new_n739), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n510), .B1(new_n776), .B2(new_n738), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n798), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n800), .A2(new_n632), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT121), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT57), .B1(new_n768), .B2(new_n510), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n838), .A4(new_n841), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(G148gat), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n833), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n632), .A2(G148gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n824), .A2(new_n481), .A3(new_n825), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT122), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n846), .A2(G148gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n848), .B1(new_n856), .B2(new_n843), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(new_n852), .C1(new_n857), .C2(new_n833), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n858), .ZN(G1345gat));
  OAI21_X1  g658(.A(G155gat), .B1(new_n817), .B2(new_n775), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n541), .A2(new_n259), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n826), .B2(new_n861), .ZN(G1346gat));
  NOR3_X1   g661(.A1(new_n817), .A2(new_n260), .A3(new_n575), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n826), .A2(new_n575), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n260), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n768), .A2(new_n319), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n601), .A3(new_n475), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT123), .ZN(new_n868));
  AOI21_X1  g667(.A(G169gat), .B1(new_n868), .B2(new_n244), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n601), .A2(new_n598), .A3(new_n468), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT124), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n779), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n244), .A2(G169gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(G1348gat));
  INV_X1    g674(.A(G176gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n876), .A3(new_n595), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n595), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(new_n876), .ZN(G1349gat));
  NAND3_X1  g679(.A1(new_n779), .A2(new_n626), .A3(new_n872), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G183gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n541), .A2(new_n347), .A3(new_n349), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n867), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT60), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n352), .A3(new_n630), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n779), .A2(new_n630), .A3(new_n872), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(G190gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n352), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n892), .A2(new_n895), .B1(new_n891), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n890), .B1(new_n894), .B2(new_n896), .ZN(G1351gat));
  AND3_X1   g696(.A1(new_n866), .A2(new_n601), .A3(new_n821), .ZN(new_n898));
  AOI21_X1  g697(.A(G197gat), .B1(new_n898), .B2(new_n244), .ZN(new_n899));
  INV_X1    g698(.A(new_n840), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n601), .A2(new_n517), .A3(new_n598), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT126), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n244), .A2(G197gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(G1352gat));
  INV_X1    g705(.A(G204gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n898), .A2(new_n907), .A3(new_n595), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT62), .Z(new_n909));
  OAI21_X1  g708(.A(G204gat), .B1(new_n903), .B2(new_n632), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1353gat));
  NAND2_X1  g710(.A1(new_n904), .A2(new_n541), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G211gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT63), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n915), .A3(G211gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n331), .A3(new_n541), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT127), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n916), .A3(new_n918), .ZN(G1354gat));
  OAI21_X1  g718(.A(G218gat), .B1(new_n903), .B2(new_n575), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n332), .A3(new_n630), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1355gat));
endmodule


