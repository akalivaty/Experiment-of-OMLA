//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n203), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n234), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT68), .A2(G1), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n253), .A2(G13), .A3(G20), .A4(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT68), .A2(G1), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT68), .A2(G1), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n257), .A2(new_n258), .A3(new_n213), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n212), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(G50), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n213), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n213), .A2(new_n267), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n264), .A2(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT72), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n272), .B1(new_n266), .B2(new_n268), .C1(new_n264), .C2(new_n265), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n261), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n212), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G41), .A2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n252), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n281), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n253), .A2(new_n254), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT69), .B1(new_n289), .B2(new_n283), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n257), .A2(new_n258), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(new_n284), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n286), .B1(new_n294), .B2(G226), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  AND4_X1   g0102(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(KEYINPUT71), .A3(G222), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n302), .ZN(new_n306));
  INV_X1    g0106(.A(G222), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(G223), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n310), .A2(new_n222), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(G190), .B(new_n295), .C1(new_n316), .C2(new_n287), .ZN(new_n317));
  INV_X1    g0117(.A(new_n295), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n287), .B1(new_n309), .B2(new_n315), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n320), .A3(KEYINPUT75), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT10), .B1(new_n278), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n276), .B(KEYINPUT9), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n318), .A2(new_n319), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(G190), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT10), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n323), .A2(new_n326), .A3(new_n327), .A4(new_n320), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n318), .B2(new_n319), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n276), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n255), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n222), .ZN(new_n337));
  INV_X1    g0137(.A(new_n262), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n222), .ZN(new_n339));
  INV_X1    g0139(.A(new_n264), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G20), .A2(G33), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G20), .B2(G77), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT74), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n265), .ZN(new_n345));
  INV_X1    g0145(.A(new_n344), .ZN(new_n346));
  INV_X1    g0146(.A(new_n265), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(KEYINPUT74), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n342), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n339), .B1(new_n261), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(KEYINPUT73), .A2(G107), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT73), .A2(G107), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n296), .A2(new_n298), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n355), .B1(new_n306), .B2(new_n236), .C1(new_n217), .C2(new_n311), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n288), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n294), .A2(G244), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n285), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n350), .B1(new_n359), .B2(new_n332), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n286), .B1(new_n356), .B2(new_n288), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n330), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n350), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n361), .B2(new_n358), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n335), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n255), .A2(G68), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT12), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n371), .B(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n202), .B2(new_n338), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n265), .A2(new_n222), .B1(new_n213), .B2(G68), .ZN(new_n375));
  INV_X1    g0175(.A(G50), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n268), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n261), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g0178(.A(new_n378), .B(KEYINPUT11), .Z(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n290), .A2(new_n293), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(G238), .A3(new_n287), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n300), .A2(new_n302), .A3(G226), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G232), .A2(G1698), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n354), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G97), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n267), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n288), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(new_n285), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n286), .B1(new_n294), .B2(G238), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n390), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n382), .B(G169), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n393), .A3(new_n390), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(G179), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n382), .B1(new_n401), .B2(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n381), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n392), .B2(new_n395), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n398), .A3(G190), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n380), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n329), .A2(new_n370), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  MUX2_X1   g0207(.A(new_n336), .B(new_n262), .S(new_n340), .Z(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT81), .Z(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT76), .B(new_n410), .C1(new_n310), .C2(G20), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(G20), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n354), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n297), .A2(G33), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n213), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT76), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G58), .A2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n213), .B1(new_n203), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n341), .A2(G159), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n421), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G58), .A2(G68), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n423), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  AOI21_X1  g0235(.A(G20), .B1(new_n296), .B2(new_n298), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(KEYINPUT7), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n413), .A3(new_n411), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n430), .B1(new_n438), .B2(G68), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(KEYINPUT78), .A3(KEYINPUT16), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n275), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n415), .A2(KEYINPUT79), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n412), .C1(new_n354), .C2(KEYINPUT79), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n410), .B1(new_n310), .B2(G20), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n202), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n431), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n442), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n409), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n286), .B1(new_n294), .B2(G232), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n310), .A2(G226), .A3(G1698), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n453), .B1(new_n267), .B2(new_n218), .C1(new_n312), .C2(new_n306), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n288), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n330), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(G169), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT18), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n432), .A2(new_n433), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT78), .B1(new_n439), .B2(KEYINPUT16), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n450), .B(new_n261), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n409), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n458), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n456), .A2(new_n367), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G190), .B2(new_n456), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n462), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT17), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n462), .A2(KEYINPUT17), .A3(new_n463), .A4(new_n469), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n459), .A2(new_n467), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n407), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT91), .B(KEYINPUT22), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n310), .A2(new_n476), .A3(new_n213), .A4(G87), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n296), .A2(new_n298), .A3(new_n213), .A4(G87), .ZN(new_n478));
  XOR2_X1   g0278(.A(KEYINPUT91), .B(KEYINPUT22), .Z(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n224), .A3(G20), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n265), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n351), .A2(G20), .A3(new_n352), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT23), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n477), .A2(new_n480), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(KEYINPUT23), .B2(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(new_n477), .A4(new_n480), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n261), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n255), .A2(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT25), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n253), .A2(G33), .A3(new_n254), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n255), .A2(new_n275), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT92), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n275), .B1(new_n489), .B2(new_n492), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT92), .B1(new_n504), .B2(new_n500), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n310), .A2(G257), .A3(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n219), .C2(new_n306), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n288), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n253), .A2(G45), .A3(new_n254), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT5), .B(G41), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n288), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G264), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n282), .A2(new_n291), .A3(new_n512), .A4(G45), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G169), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n508), .A2(new_n288), .B1(new_n513), .B2(G264), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G179), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n503), .A2(new_n505), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n509), .A2(new_n514), .A3(new_n365), .A4(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT93), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n518), .A2(new_n524), .A3(new_n365), .A4(new_n515), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n516), .A2(new_n367), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n504), .A2(new_n500), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g0330(.A(KEYINPUT73), .B(G107), .Z(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n444), .B2(new_n445), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  XNOR2_X1  g0333(.A(G97), .B(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n213), .B1(new_n222), .B2(new_n268), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n261), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT82), .B1(new_n255), .B2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n336), .A2(new_n540), .A3(new_n388), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n539), .A2(new_n541), .B1(new_n498), .B2(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT83), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n303), .A2(KEYINPUT84), .A3(KEYINPUT4), .A4(G244), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT70), .B(G1698), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n310), .A2(new_n548), .A3(KEYINPUT4), .A4(G244), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n306), .B2(new_n223), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(G1698), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n547), .A2(new_n551), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n288), .ZN(new_n558));
  AND2_X1   g0358(.A1(KEYINPUT5), .A2(G41), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT5), .A2(G41), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(new_n287), .C1(new_n510), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n515), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G200), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  AOI211_X1 g0365(.A(G190), .B(new_n563), .C1(new_n557), .C2(new_n288), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n545), .B(new_n546), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n332), .B1(new_n558), .B2(new_n564), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n330), .B(new_n563), .C1(new_n557), .C2(new_n288), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n543), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G87), .A2(G97), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n531), .A2(new_n571), .B1(new_n213), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n296), .A2(new_n298), .A3(new_n213), .A4(G68), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n265), .B2(new_n388), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n261), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n336), .A2(new_n344), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n498), .A2(new_n346), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n296), .A2(new_n298), .A3(G244), .A4(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G116), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n306), .C2(new_n217), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n310), .A2(new_n548), .A3(G238), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n583), .A4(new_n584), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n288), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n510), .A2(new_n219), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n291), .A2(G45), .A3(new_n279), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n287), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n330), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n593), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n287), .B1(new_n585), .B2(KEYINPUT85), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n589), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n582), .B(new_n594), .C1(G169), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n590), .A2(G190), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n498), .A2(G87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n578), .A2(new_n579), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n599), .B(new_n602), .C1(new_n367), .C2(new_n597), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n567), .A2(new_n570), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n530), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n558), .A2(new_n564), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n563), .B1(new_n557), .B2(new_n288), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G179), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n558), .A2(new_n365), .A3(new_n564), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G200), .B2(new_n609), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT83), .B1(new_n538), .B2(new_n542), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n543), .A2(new_n611), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n590), .A2(new_n593), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n332), .B1(new_n580), .B2(new_n581), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n601), .B1(new_n597), .B2(G190), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(G200), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n619), .A2(new_n594), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(KEYINPUT86), .A3(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n260), .A2(new_n212), .B1(G20), .B2(new_n483), .ZN(new_n624));
  AOI21_X1  g0424(.A(G20), .B1(G33), .B2(G283), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n267), .A2(G97), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n625), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(KEYINPUT20), .B(new_n624), .C1(new_n628), .C2(new_n629), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(KEYINPUT90), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n255), .A2(new_n483), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n498), .B2(new_n483), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n637), .A3(new_n631), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n296), .A2(new_n298), .A3(G257), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n300), .A2(new_n302), .ZN(new_n641));
  AND2_X1   g0441(.A1(KEYINPUT87), .A2(G303), .ZN(new_n642));
  NOR2_X1   g0442(.A1(KEYINPUT87), .A2(G303), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n640), .A2(new_n641), .B1(new_n644), .B2(new_n310), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n310), .A2(G264), .A3(G1698), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n288), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(KEYINPUT88), .B(new_n288), .C1(new_n645), .C2(new_n647), .ZN(new_n651));
  OAI211_X1 g0451(.A(G270), .B(new_n287), .C1(new_n510), .C2(new_n561), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n515), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n639), .B1(G200), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n365), .B2(new_n654), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT21), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n653), .ZN(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT87), .B(G303), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n354), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n646), .B(new_n660), .C1(new_n641), .C2(new_n640), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT88), .B1(new_n661), .B2(new_n288), .ZN(new_n662));
  OAI21_X1  g0462(.A(G169), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n633), .A2(KEYINPUT90), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n625), .A2(new_n626), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT89), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT20), .B1(new_n668), .B2(new_n624), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n636), .A2(new_n638), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n657), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n658), .A2(new_n662), .A3(new_n330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n639), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n654), .A2(new_n639), .A3(KEYINPUT21), .A4(G169), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n656), .A2(new_n673), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n475), .A2(new_n606), .A3(new_n623), .A4(new_n678), .ZN(G372));
  INV_X1    g0479(.A(new_n403), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n406), .B2(new_n364), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n472), .A2(new_n473), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n459), .B(new_n467), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n329), .B(KEYINPUT94), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n335), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n622), .A2(new_n529), .A3(new_n570), .A4(new_n567), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n516), .A2(new_n330), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n332), .B1(new_n518), .B2(new_n515), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n504), .B2(new_n500), .ZN(new_n689));
  AND4_X1   g0489(.A1(new_n673), .A2(new_n689), .A3(new_n675), .A4(new_n676), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  INV_X1    g0492(.A(new_n616), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n622), .A2(new_n692), .A3(new_n611), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n598), .A2(new_n603), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT26), .B1(new_n695), .B2(new_n570), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n696), .A3(new_n598), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n475), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n685), .A2(new_n698), .ZN(G369));
  AND2_X1   g0499(.A1(new_n213), .A2(G13), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n291), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  OAI21_X1  g0502(.A(G213), .B1(new_n701), .B2(KEYINPUT27), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n639), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT95), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n677), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT96), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n677), .A2(new_n709), .ZN(new_n715));
  INV_X1    g0515(.A(new_n713), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT96), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n503), .A2(new_n505), .A3(new_n707), .ZN(new_n718));
  INV_X1    g0518(.A(new_n707), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n530), .A2(new_n718), .B1(new_n521), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n714), .A2(new_n717), .A3(new_n720), .A4(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n689), .A2(new_n707), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n712), .A2(new_n719), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n530), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n207), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G1), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n531), .A2(new_n483), .A3(new_n571), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(new_n210), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n719), .B1(new_n697), .B2(new_n691), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT97), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n719), .C1(new_n697), .C2(new_n691), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n503), .A2(new_n505), .A3(new_n520), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n712), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n686), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n568), .A2(new_n569), .B1(new_n614), .B2(new_n615), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT26), .B1(new_n695), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n543), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n608), .B2(new_n610), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n692), .A3(new_n598), .A4(new_n603), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n748), .A3(new_n598), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT29), .B(new_n719), .C1(new_n743), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n521), .A2(new_n673), .A3(new_n675), .A4(new_n676), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n617), .A3(new_n529), .A4(new_n622), .ZN(new_n754));
  INV_X1    g0554(.A(new_n598), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n695), .A2(new_n570), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n692), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n745), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(KEYINPUT98), .A3(KEYINPUT29), .A4(new_n719), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n740), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n606), .A2(new_n623), .A3(new_n678), .A4(new_n719), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n674), .A2(new_n518), .A3(new_n609), .A4(new_n597), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n609), .A2(new_n518), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(KEYINPUT30), .A3(new_n597), .A4(new_n674), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n654), .A2(new_n618), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n516), .A2(new_n330), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n609), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n765), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n707), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT31), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n763), .A2(new_n764), .B1(new_n770), .B2(new_n768), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n719), .B1(new_n776), .B2(new_n767), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT31), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n762), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G330), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n761), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT99), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n761), .A2(KEYINPUT99), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n734), .B1(new_n785), .B2(G1), .ZN(G364));
  NAND3_X1  g0586(.A1(new_n714), .A2(new_n717), .A3(G330), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n252), .B1(new_n700), .B2(G45), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n729), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(G330), .B1(new_n714), .B2(new_n717), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n710), .A2(new_n713), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n728), .A2(new_n354), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G355), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G116), .B2(new_n207), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n249), .A2(G45), .ZN(new_n802));
  INV_X1    g0602(.A(G45), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n310), .B(new_n728), .C1(new_n211), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n212), .B1(G20), .B2(new_n332), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT100), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n790), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n213), .A2(new_n330), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n811), .A2(new_n367), .A3(G190), .ZN(new_n812));
  NOR2_X1   g0612(.A1(KEYINPUT33), .A2(G317), .ZN(new_n813));
  AND2_X1   g0613(.A1(KEYINPUT33), .A2(G317), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G190), .A2(G200), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n365), .A2(new_n367), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n810), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(G326), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n365), .A2(G179), .A3(G200), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n213), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G294), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n811), .A2(new_n365), .A3(G200), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n213), .A2(G179), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n817), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n828), .A2(G322), .B1(G329), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n820), .A2(new_n829), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n310), .B1(new_n834), .B2(G303), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n829), .A2(new_n365), .A3(G200), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT103), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G283), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n823), .A2(new_n827), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(G107), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n310), .B1(new_n833), .B2(new_n218), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT104), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n830), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G97), .B2(new_n826), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n828), .A2(G58), .B1(new_n822), .B2(G50), .ZN(new_n852));
  INV_X1    g0652(.A(new_n818), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n812), .A2(G68), .B1(G77), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n840), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n809), .B1(new_n856), .B2(new_n806), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n792), .A2(new_n794), .B1(new_n798), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G396));
  OAI22_X1  g0659(.A1(new_n366), .A2(new_n368), .B1(new_n350), .B2(new_n719), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n363), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT108), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n360), .A2(new_n362), .A3(new_n719), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(KEYINPUT109), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT109), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n736), .A3(new_n739), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n694), .A2(new_n598), .A3(new_n696), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n686), .A2(new_n690), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n707), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n790), .B1(new_n876), .B2(new_n780), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n780), .B2(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(new_n806), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n812), .A2(G150), .B1(new_n822), .B2(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  INV_X1    g0681(.A(new_n828), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .C1(new_n847), .C2(new_n818), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n838), .A2(G68), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n310), .B1(new_n830), .B2(new_n886), .C1(new_n376), .C2(new_n833), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G58), .B2(new_n826), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n812), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(G283), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n893), .A2(new_n894), .B1(new_n483), .B2(new_n818), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT106), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n838), .A2(G87), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n354), .B1(new_n833), .B2(new_n224), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n828), .A2(G294), .B1(new_n822), .B2(G303), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n816), .B2(new_n830), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n898), .B(new_n900), .C1(G97), .C2(new_n826), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n895), .A2(KEYINPUT106), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n889), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n879), .B1(new_n904), .B2(KEYINPUT107), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(KEYINPUT107), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n806), .A2(new_n795), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n791), .B1(new_n222), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n906), .B(new_n908), .C1(new_n796), .C2(new_n866), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n878), .A2(new_n909), .ZN(G384));
  INV_X1    g0710(.A(new_n536), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n214), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  NAND3_X1  g0715(.A1(new_n211), .A2(G77), .A3(new_n421), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n376), .A2(G68), .ZN(new_n917));
  AOI211_X1 g0717(.A(G13), .B(new_n291), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n863), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n874), .B2(new_n866), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT110), .ZN(new_n923));
  OAI21_X1  g0723(.A(G169), .B1(new_n392), .B2(new_n395), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT14), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n406), .A2(new_n925), .A3(new_n399), .A4(new_n396), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n380), .A2(new_n719), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n403), .A2(new_n406), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n926), .A2(new_n923), .A3(new_n927), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n439), .A2(KEYINPUT16), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n408), .B1(new_n441), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n470), .B1(new_n935), .B2(new_n705), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n458), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n464), .A2(new_n465), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n464), .A2(new_n704), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT37), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n470), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n935), .A2(new_n705), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n474), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n943), .A2(new_n945), .A3(KEYINPUT38), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n922), .B(new_n933), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n459), .A2(new_n467), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n705), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n680), .A2(new_n719), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n470), .B1(new_n451), .B2(new_n458), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n451), .A2(new_n705), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT37), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT111), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(new_n942), .ZN(new_n958));
  OAI211_X1 g0758(.A(KEYINPUT111), .B(KEYINPUT37), .C1(new_n954), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n474), .A2(new_n955), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT38), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n942), .A2(new_n938), .B1(new_n474), .B2(new_n944), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT39), .B1(new_n964), .B2(KEYINPUT38), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT39), .B1(new_n947), .B2(new_n946), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n951), .B1(new_n953), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n740), .A2(new_n760), .A3(new_n475), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n685), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n931), .A2(new_n866), .A3(new_n932), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n774), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n777), .B2(KEYINPUT31), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n762), .A2(new_n778), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n973), .B(new_n977), .C1(new_n947), .C2(new_n946), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT40), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n964), .A2(KEYINPUT38), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n963), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n973), .A2(KEYINPUT40), .A3(new_n977), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n984), .A3(new_n475), .A4(new_n977), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(G330), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n980), .A2(new_n984), .B1(new_n475), .B2(new_n977), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n972), .A2(new_n988), .B1(new_n291), .B2(new_n700), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n972), .A2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n919), .B1(new_n989), .B2(new_n990), .ZN(G367));
  NOR2_X1   g0791(.A1(new_n728), .A2(new_n310), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n234), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n808), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n207), .B2(new_n344), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n790), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n882), .A2(new_n644), .B1(new_n821), .B2(new_n816), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n818), .A2(new_n894), .B1(new_n830), .B2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n354), .B1(new_n837), .B2(new_n388), .C1(new_n825), .C2(new_n531), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n834), .A2(G116), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT46), .ZN(new_n1003));
  INV_X1    g0803(.A(G294), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1001), .B(new_n1003), .C1(new_n1004), .C2(new_n893), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n826), .A2(G68), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n881), .B2(new_n821), .C1(new_n882), .C2(new_n266), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT118), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n310), .B1(new_n837), .B2(new_n222), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n833), .A2(new_n201), .B1(new_n830), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G50), .C2(new_n853), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n893), .B2(new_n847), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1005), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n996), .B1(new_n1015), .B2(new_n806), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n622), .B1(new_n602), .B2(new_n719), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n755), .A2(new_n601), .A3(new_n707), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n1018), .A3(new_n797), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT116), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n707), .B1(new_n614), .B2(new_n615), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n567), .A2(new_n570), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT114), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT114), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n567), .A2(new_n570), .A3(new_n1025), .A4(new_n1022), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n744), .A2(new_n719), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n726), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1031), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n725), .ZN(new_n1035));
  AND4_X1   g0835(.A1(KEYINPUT44), .A2(new_n1027), .A3(new_n725), .A4(new_n1029), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT44), .B1(new_n1034), .B2(new_n725), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1032), .B(new_n1035), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n721), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1027), .A2(new_n725), .A3(new_n1029), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT44), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1034), .A2(KEYINPUT44), .A3(new_n725), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1045), .A2(new_n721), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n724), .A2(new_n530), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n724), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n720), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n787), .B(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n783), .A2(new_n784), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n729), .B(KEYINPUT41), .Z(new_n1055));
  OAI21_X1  g0855(.A(new_n1021), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI221_X4 g0856(.A(new_n782), .B1(G330), .B2(new_n779), .C1(new_n740), .C2(new_n760), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT99), .B1(new_n761), .B2(new_n780), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1057), .A2(new_n1058), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1055), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(KEYINPUT116), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n789), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT117), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1030), .A2(new_n1048), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT42), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n570), .B1(new_n1034), .B2(new_n521), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n719), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n1071), .A2(KEYINPUT43), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1069), .A2(KEYINPUT43), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n721), .A2(new_n1034), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1075), .B(new_n1079), .C1(new_n1068), .C2(new_n1077), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1063), .A2(new_n1064), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1060), .A2(KEYINPUT116), .A3(new_n1061), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT116), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n788), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT117), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1020), .B1(new_n1084), .B2(new_n1089), .ZN(G387));
  AOI21_X1  g0890(.A(new_n1052), .B1(new_n783), .B2(new_n784), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n730), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n785), .B2(new_n1053), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1053), .A2(new_n789), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n797), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n720), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n354), .B1(new_n837), .B2(new_n483), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT121), .B(G322), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n822), .A2(new_n1099), .B1(new_n853), .B2(new_n659), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n998), .B2(new_n882), .C1(new_n893), .C2(new_n816), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n826), .A2(G283), .B1(new_n834), .B2(G294), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT49), .Z(new_n1107));
  AOI211_X1 g0907(.A(new_n1097), .B(new_n1107), .C1(G326), .C2(new_n831), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n828), .A2(G50), .B1(G150), .B2(new_n831), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n847), .B2(new_n821), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n812), .A2(new_n340), .B1(G68), .B2(new_n853), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n826), .A2(new_n346), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n834), .A2(G77), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n310), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1110), .B(new_n1114), .C1(G97), .C2(new_n838), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n806), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n732), .A2(new_n799), .B1(new_n224), .B2(new_n728), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n732), .B(KEYINPUT119), .Z(new_n1118));
  OAI21_X1  g0918(.A(new_n803), .B1(new_n202), .B2(new_n222), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n264), .A2(G50), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT50), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n992), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1124), .A2(KEYINPUT120), .B1(new_n803), .B2(new_n239), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(KEYINPUT120), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1117), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n791), .B1(new_n1127), .B2(new_n994), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1093), .B(new_n1094), .C1(new_n1096), .C2(new_n1129), .ZN(G393));
  NAND2_X1  g0930(.A1(new_n1047), .A2(new_n789), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n245), .A2(new_n992), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n808), .B1(G97), .B2(new_n728), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n791), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n893), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n659), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n828), .A2(G311), .B1(new_n822), .B2(G317), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT52), .Z(new_n1138));
  OAI21_X1  g0938(.A(new_n354), .B1(new_n818), .B2(new_n1004), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n833), .A2(new_n894), .B1(new_n830), .B2(new_n1098), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G116), .C2(new_n826), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1136), .A2(new_n841), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1135), .A2(G50), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n828), .A2(G159), .B1(new_n822), .B2(G150), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT51), .Z(new_n1145));
  OAI22_X1  g0945(.A1(new_n818), .A2(new_n264), .B1(new_n830), .B2(new_n881), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n825), .A2(new_n222), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n310), .B1(new_n833), .B2(new_n202), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1143), .A2(new_n897), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1142), .A2(new_n1150), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1134), .B1(new_n879), .B2(new_n1151), .C1(new_n1030), .C2(new_n1095), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1131), .A2(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1091), .A2(new_n1047), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n730), .B1(new_n1091), .B2(new_n1047), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G390));
  NAND2_X1  g0957(.A1(new_n931), .A2(new_n932), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n952), .B1(new_n921), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n966), .A2(new_n1159), .A3(new_n967), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n758), .A2(new_n866), .A3(new_n719), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n863), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n953), .B1(new_n1162), .B2(new_n933), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n982), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n973), .A2(G330), .A3(new_n977), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n977), .A2(new_n475), .A3(G330), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n970), .A2(new_n685), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n779), .A2(G330), .A3(new_n866), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n1158), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n922), .B1(new_n1172), .B2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n977), .A2(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1158), .B1(new_n1174), .B2(new_n870), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1162), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n933), .A2(new_n779), .A3(G330), .A4(new_n866), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1170), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1160), .A2(new_n1164), .A3(new_n1177), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1168), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1181), .A2(new_n729), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n1170), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1168), .A2(new_n1180), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(KEYINPUT122), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1186), .A2(new_n788), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1135), .A2(new_n353), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n821), .A2(new_n894), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n818), .A2(new_n388), .B1(new_n830), .B2(new_n1004), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G116), .C2(new_n828), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n310), .B(new_n1147), .C1(G87), .C2(new_n834), .ZN(new_n1195));
  AND4_X1   g0995(.A1(new_n885), .A2(new_n1191), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n833), .A2(new_n266), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT53), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n893), .B2(new_n1010), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT54), .B(G143), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n882), .A2(new_n886), .B1(new_n818), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(G128), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1202), .A2(new_n821), .B1(new_n837), .B2(new_n376), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n354), .B1(new_n831), .B2(G125), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n847), .B2(new_n825), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1199), .A2(new_n1201), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n806), .B1(new_n1196), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n907), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n790), .C1(new_n340), .C2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n966), .A2(new_n967), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n795), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1190), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1189), .A2(new_n1212), .ZN(G378));
  INV_X1    g1013(.A(G330), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n978), .B2(new_n979), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n984), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n276), .A2(new_n704), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT55), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n684), .A2(new_n334), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n684), .B2(new_n334), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1218), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n684), .A2(new_n334), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1220), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n684), .A2(new_n334), .A3(new_n1221), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1217), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1216), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1215), .A2(new_n984), .A3(new_n1229), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n969), .A3(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n948), .B(new_n950), .C1(new_n1210), .C2(new_n952), .ZN(new_n1234));
  AND4_X1   g1034(.A1(G330), .A2(new_n980), .A3(new_n984), .A4(new_n1229), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1229), .B1(new_n1215), .B2(new_n984), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1170), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1233), .A2(new_n1237), .B1(new_n1181), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n729), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1181), .A2(new_n1238), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1241), .A2(KEYINPUT57), .A3(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n791), .B1(new_n376), .B2(new_n907), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n890), .A2(new_n886), .B1(new_n833), .B2(new_n1200), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n828), .A2(G128), .B1(new_n822), .B2(G125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1010), .B2(new_n818), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G150), .C2(new_n826), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G33), .A2(G41), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT123), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n837), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1256), .A2(G159), .B1(new_n831), .B2(G124), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1251), .A2(new_n1252), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n812), .A2(G97), .B1(G58), .B2(new_n1256), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n310), .A2(G41), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n1006), .A3(new_n1113), .A4(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n818), .A2(new_n344), .B1(new_n830), .B2(new_n894), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n882), .A2(new_n224), .B1(new_n821), .B2(new_n483), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT58), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1254), .B(new_n376), .C1(G41), .C2(new_n310), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1264), .A2(KEYINPUT58), .ZN(new_n1267));
  AND4_X1   g1067(.A1(new_n1258), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1245), .B1(new_n879), .B2(new_n1268), .C1(new_n1229), .C2(new_n796), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT125), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(KEYINPUT125), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1241), .A2(new_n789), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1244), .A2(new_n1272), .ZN(G375));
  AND3_X1   g1073(.A1(new_n1173), .A2(new_n1170), .A3(new_n1178), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1185), .A2(new_n1061), .A3(new_n1187), .A4(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n791), .B1(new_n202), .B2(new_n907), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n893), .A2(new_n1200), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G159), .A2(new_n834), .B1(new_n831), .B2(G128), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n266), .B2(new_n818), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n828), .A2(G137), .B1(new_n822), .B2(G132), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n376), .B2(new_n825), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1278), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n310), .B1(new_n837), .B2(new_n201), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT126), .Z(new_n1285));
  AOI22_X1  g1085(.A1(new_n1135), .A2(G116), .B1(G77), .B2(new_n838), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n353), .A2(new_n853), .B1(new_n831), .B2(G303), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1287), .B1(new_n1004), .B2(new_n821), .C1(new_n894), .C2(new_n882), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1112), .B(new_n354), .C1(new_n388), .C2(new_n833), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1283), .A2(new_n1285), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1277), .B1(new_n879), .B2(new_n1291), .C1(new_n933), .C2(new_n796), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1184), .B2(new_n788), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1276), .A2(new_n1294), .ZN(G381));
  INV_X1    g1095(.A(G384), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1156), .A2(new_n1296), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G393), .A2(new_n1297), .A3(G381), .A4(G396), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1211), .B(new_n1190), .C1(new_n1182), .C2(new_n1188), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OR3_X1    g1100(.A1(G375), .A2(new_n1300), .A3(G387), .ZN(G407));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n706), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G407), .B(G213), .C1(G375), .C2(new_n1302), .ZN(G409));
  OAI21_X1  g1103(.A(new_n1064), .B1(new_n1063), .B2(new_n1083), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n1088), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G390), .B1(new_n1306), .B2(new_n1020), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1020), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1308), .B(new_n1156), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(G396), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(new_n858), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G387), .A2(new_n1156), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1306), .A2(new_n1020), .A3(G390), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G378), .B(new_n1272), .C1(new_n1240), .C2(new_n1243), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1241), .A2(new_n1061), .A3(new_n1242), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1272), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1299), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(G213), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(G343), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT60), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1179), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n730), .B1(new_n1329), .B2(new_n1274), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1275), .B1(new_n1328), .B2(new_n1179), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G384), .B1(new_n1332), .B2(new_n1294), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1293), .B(new_n1296), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1327), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1329), .A2(new_n1274), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1184), .A2(KEYINPUT60), .A3(new_n1170), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n729), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1296), .B1(new_n1339), .B2(new_n1293), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1332), .A2(G384), .A3(new_n1294), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1341), .A3(new_n1326), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1335), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1323), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(KEYINPUT63), .A3(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1321), .A2(new_n1348), .A3(new_n1324), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1316), .A2(new_n1345), .A3(new_n1349), .A4(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1346), .B2(new_n1343), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT62), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1350), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1346), .A2(KEYINPUT62), .A3(new_n1348), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1355), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1353), .B1(new_n1316), .B2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1299), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1347), .A2(KEYINPUT127), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1363), .A3(new_n1317), .ZN(new_n1364));
  AOI21_X1  g1164(.A(G378), .B1(new_n1244), .B2(new_n1272), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1317), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1362), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1364), .A2(new_n1367), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1316), .A2(new_n1364), .A3(new_n1367), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(G402));
endmodule


