//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  AOI22_X1  g053(.A1(G124), .A2(new_n477), .B1(new_n478), .B2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  INV_X1    g055(.A(new_n469), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n472), .A2(KEYINPUT70), .A3(G138), .A4(new_n462), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G102), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n501), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  INV_X1    g089(.A(G51), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(G89), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n505), .A2(new_n515), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G168));
  NAND2_X1  g097(.A1(G77), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  INV_X1    g099(.A(G64), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n511), .B1(new_n526), .B2(KEYINPUT72), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n527), .B1(KEYINPUT72), .B2(new_n526), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n502), .A2(new_n503), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G52), .Z(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G90), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n537), .A2(new_n505), .B1(new_n507), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  XOR2_X1   g121(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n547));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n532), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n524), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  NAND2_X1  g133(.A1(new_n530), .A2(G87), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n532), .A2(G49), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G288));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n507), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n530), .A2(KEYINPUT76), .A3(G86), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n532), .B2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n511), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n530), .A2(G85), .B1(new_n532), .B2(G47), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT77), .ZN(G290));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  OR3_X1    g158(.A1(G171), .A2(KEYINPUT78), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n530), .A2(G92), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT10), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G54), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n511), .A2(new_n587), .B1(new_n505), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT78), .B1(new_n591), .B2(new_n583), .ZN(new_n592));
  NOR2_X1   g167(.A1(G171), .A2(new_n583), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n592), .B2(new_n593), .ZN(G284));
  OAI21_X1  g169(.A(new_n584), .B1(new_n592), .B2(new_n593), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(KEYINPUT79), .B1(G299), .B2(new_n583), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT79), .B2(new_n596), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(KEYINPUT79), .B2(new_n596), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(G860), .ZN(G148));
  NOR2_X1   g176(.A1(new_n542), .A2(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n591), .A2(G559), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n469), .A2(G2104), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n469), .A2(G135), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT80), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n477), .A2(G123), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT81), .ZN(new_n613));
  AND2_X1   g188(.A1(G111), .A2(G2105), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G99), .B2(new_n462), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n611), .B(new_n613), .C1(new_n466), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XOR2_X1   g196(.A(G2443), .B(G2446), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT84), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n628), .B2(new_n630), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(G401));
  XNOR2_X1  g210(.A(G2072), .B(G2078), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT85), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2084), .B(G2090), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n643));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n644), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n641), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  OR3_X1    g236(.A1(new_n652), .A2(new_n655), .A3(new_n660), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G229));
  NAND2_X1  g244(.A1(new_n477), .A2(G129), .ZN(new_n670));
  NAND3_X1  g245(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n469), .A2(G141), .ZN(new_n675));
  AND4_X1   g250(.A1(new_n670), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(G32), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT27), .B(G1996), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT99), .Z(new_n682));
  AND2_X1   g257(.A1(KEYINPUT24), .A2(G34), .ZN(new_n683));
  NOR2_X1   g258(.A1(KEYINPUT24), .A2(G34), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n677), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G160), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n677), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n682), .B1(G2084), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G29), .A2(G33), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n469), .A2(G139), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT25), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(KEYINPUT25), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n472), .A2(G127), .ZN(new_n698));
  INV_X1    g273(.A(G115), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n466), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n462), .B1(new_n700), .B2(KEYINPUT96), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(KEYINPUT96), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n690), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G2072), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT31), .B(G11), .Z(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT101), .Z(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n716), .B2(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n714), .B(new_n720), .C1(new_n677), .C2(new_n616), .ZN(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G171), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT102), .Z(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n724), .B2(G1961), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT103), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G35), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G162), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n710), .A2(G20), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT105), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT23), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G299), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1956), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n677), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n477), .A2(G128), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT92), .ZN(new_n743));
  MUX2_X1   g318(.A(G104), .B(G116), .S(G2105), .Z(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(G2104), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n469), .A2(G140), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT91), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G164), .A2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G27), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT104), .B(G2078), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n738), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n724), .A2(G1961), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n688), .A2(G2084), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n757), .B1(new_n753), .B2(new_n754), .C1(new_n679), .C2(new_n680), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n543), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n590), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1348), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n758), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n732), .A2(new_n755), .A3(new_n756), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n709), .A2(new_n726), .A3(new_n727), .A4(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n710), .A2(G23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n563), .B2(new_n710), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT33), .B(G1976), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G22), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT89), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G303), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1971), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n770), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(KEYINPUT34), .ZN(new_n780));
  AOI22_X1  g355(.A1(G119), .A2(new_n477), .B1(new_n469), .B2(G131), .ZN(new_n781));
  INV_X1    g356(.A(G95), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(new_n462), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT87), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT88), .Z(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  XOR2_X1   g363(.A(KEYINPUT35), .B(G1991), .Z(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(G16), .A2(G24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G290), .B2(new_n710), .ZN(new_n793));
  INV_X1    g368(.A(G1986), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n780), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT90), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n779), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT36), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n797), .A2(new_n801), .A3(new_n798), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n767), .B1(new_n800), .B2(new_n802), .ZN(G311));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n802), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n709), .A2(new_n726), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n804), .A2(new_n727), .A3(new_n766), .A4(new_n805), .ZN(G150));
  NAND2_X1  g381(.A1(new_n590), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n542), .A2(KEYINPUT106), .ZN(new_n809));
  INV_X1    g384(.A(G55), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n810), .A2(new_n505), .B1(new_n507), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n511), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n539), .A2(KEYINPUT106), .A3(new_n541), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n809), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n815), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n818), .A2(KEYINPUT106), .A3(new_n542), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n808), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n815), .A2(new_n823), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n748), .B(new_n499), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n676), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n833), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n607), .B(new_n786), .ZN(new_n838));
  MUX2_X1   g413(.A(G106), .B(G118), .S(G2105), .Z(new_n839));
  AOI22_X1  g414(.A1(G130), .A2(new_n477), .B1(new_n839), .B2(G2104), .ZN(new_n840));
  INV_X1    g415(.A(G142), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n481), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n838), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n834), .A2(new_n843), .A3(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(new_n686), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n616), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n834), .A2(KEYINPUT108), .A3(new_n843), .A4(new_n836), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n854), .A2(new_n845), .A3(new_n855), .A4(new_n849), .ZN(new_n856));
  AND4_X1   g431(.A1(KEYINPUT40), .A2(new_n851), .A3(new_n852), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n847), .B2(new_n850), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT40), .B1(new_n858), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(G395));
  NOR2_X1   g435(.A1(new_n818), .A2(G868), .ZN(new_n861));
  XNOR2_X1  g436(.A(G290), .B(new_n562), .ZN(new_n862));
  XNOR2_X1  g437(.A(G303), .B(G305), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n590), .B(G299), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT41), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(KEYINPUT109), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n820), .B(new_n603), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n869), .B(new_n870), .S(new_n871), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n861), .B1(new_n873), .B2(G868), .ZN(G295));
  AOI21_X1  g449(.A(new_n861), .B1(new_n873), .B2(G868), .ZN(G331));
  INV_X1    g450(.A(KEYINPUT112), .ZN(new_n876));
  XNOR2_X1  g451(.A(G301), .B(G168), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n820), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n820), .A2(new_n877), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n870), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT111), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n879), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n881), .A2(new_n882), .B1(new_n869), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(KEYINPUT111), .A3(new_n870), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n864), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n868), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n869), .A2(new_n883), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n864), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n852), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n876), .B1(new_n891), .B2(KEYINPUT43), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n876), .B(KEYINPUT43), .C1(new_n886), .C2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n888), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n865), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(KEYINPUT44), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n895), .B1(new_n886), .B2(new_n890), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(KEYINPUT43), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n892), .A2(new_n899), .B1(KEYINPUT44), .B2(new_n902), .ZN(G397));
  INV_X1    g478(.A(KEYINPUT127), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n748), .A2(G2067), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT114), .ZN(new_n906));
  INV_X1    g481(.A(G2067), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n745), .B2(new_n747), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  INV_X1    g485(.A(G1996), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n909), .B(new_n910), .C1(new_n911), .C2(new_n676), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n496), .A2(new_n497), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT70), .B1(new_n469), .B2(G138), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n491), .ZN(new_n915));
  AOI21_X1  g490(.A(G1384), .B1(new_n915), .B2(new_n490), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n473), .A2(new_n474), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G2105), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(G40), .A3(new_n464), .A4(new_n470), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n916), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT113), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT113), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n923), .A3(new_n911), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n912), .A2(new_n920), .B1(new_n926), .B2(new_n676), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n786), .B(new_n790), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n920), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(new_n794), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n927), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n552), .A2(KEYINPUT57), .A3(new_n556), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n498), .A2(new_n492), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n919), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT45), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT115), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT115), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n499), .A2(new_n945), .A3(KEYINPUT45), .A4(new_n937), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT56), .B(G2072), .Z(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n942), .A2(new_n944), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n499), .A2(new_n950), .A3(new_n937), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n471), .A2(new_n475), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n499), .B2(new_n937), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n737), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n936), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n957), .A3(new_n936), .ZN(new_n959));
  INV_X1    g534(.A(G1348), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n937), .B(new_n955), .C1(new_n938), .C2(new_n939), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n953), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n950), .B1(new_n499), .B2(new_n937), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n940), .A2(new_n919), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n907), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n591), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n958), .B1(new_n959), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n949), .A2(new_n957), .A3(new_n936), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(new_n958), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT59), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n942), .A2(new_n944), .A3(new_n911), .A4(new_n946), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n916), .A2(new_n953), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT58), .B(G1341), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n971), .B1(new_n977), .B2(new_n543), .ZN(new_n978));
  AOI211_X1 g553(.A(KEYINPUT59), .B(new_n542), .C1(new_n972), .C2(new_n976), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n970), .A2(KEYINPUT61), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n949), .A2(new_n957), .ZN(new_n981));
  INV_X1    g556(.A(new_n936), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(KEYINPUT61), .A3(new_n959), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n964), .A2(new_n591), .A3(new_n966), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT60), .B1(new_n985), .B2(new_n967), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT60), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n964), .A2(new_n987), .A3(new_n590), .A4(new_n966), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n968), .B1(new_n980), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n942), .A2(new_n944), .A3(new_n991), .A4(new_n946), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  INV_X1    g568(.A(G1961), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n940), .A2(KEYINPUT50), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(new_n953), .A3(new_n961), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n953), .B1(new_n916), .B2(KEYINPUT45), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n945), .B1(new_n916), .B2(KEYINPUT45), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(KEYINPUT53), .A3(new_n991), .A4(new_n946), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1001), .A3(G301), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT124), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n997), .A2(new_n1001), .A3(KEYINPUT124), .A4(G301), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n992), .A2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n996), .A2(new_n994), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n942), .A2(KEYINPUT53), .A3(new_n991), .A4(new_n943), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G171), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1005), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1006), .A2(new_n1008), .A3(G301), .A4(new_n1007), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT54), .ZN(new_n1015));
  AOI21_X1  g590(.A(G301), .B1(new_n997), .B2(new_n1001), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n943), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n713), .B1(new_n998), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT121), .B(G2084), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n995), .A2(new_n953), .A3(new_n961), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT118), .B(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G168), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1025), .B(KEYINPUT123), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT51), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1024), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1966), .B1(new_n942), .B2(new_n943), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n962), .A2(new_n963), .A3(new_n1020), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1025), .A2(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1026), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1017), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n990), .A2(new_n1013), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT125), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1010), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n1029), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1036), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1023), .B2(new_n1032), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(KEYINPUT62), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1042), .A2(new_n1043), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1040), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n942), .A2(new_n946), .A3(new_n944), .ZN(new_n1059));
  INV_X1    g634(.A(G1971), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n954), .A2(G2090), .A3(new_n956), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT120), .B(new_n1058), .C1(new_n1063), .C2(new_n1024), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n965), .A2(new_n1024), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n563), .A2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n564), .A2(new_n1068), .A3(new_n566), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G48), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n511), .A2(new_n574), .B1(new_n505), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n507), .A2(new_n570), .ZN(new_n1073));
  OAI21_X1  g648(.A(G1981), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(G305), .B2(G1981), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1074), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1065), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n973), .A2(new_n1032), .A3(new_n1067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT52), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1070), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n996), .A2(G2090), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1027), .B1(new_n1083), .B2(new_n1061), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1084), .B2(new_n1057), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1024), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1057), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1064), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1054), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1035), .A2(G286), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1064), .A2(new_n1085), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1035), .A2(new_n1093), .A3(G286), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1085), .B(new_n1095), .C1(new_n1057), .C2(new_n1084), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1084), .A2(new_n1057), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n1082), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G305), .A2(G1981), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1079), .A2(new_n1068), .A3(new_n567), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n932), .B1(new_n1090), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT46), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n925), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n925), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n909), .A2(new_n676), .A3(new_n910), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n920), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NOR3_X1   g691(.A1(G290), .A2(new_n930), .A3(G1986), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT48), .Z(new_n1118));
  NAND3_X1  g693(.A1(new_n927), .A2(new_n929), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n787), .A2(new_n790), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n905), .B1(new_n927), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1116), .B(new_n1119), .C1(new_n930), .C2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n904), .B1(new_n1107), .B2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1121), .A2(new_n930), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1124), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1054), .B2(new_n1089), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(KEYINPUT127), .C1(new_n1127), .C2(new_n932), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g704(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n1131));
  NOR4_X1   g705(.A1(G227), .A2(new_n460), .A3(G401), .A4(G229), .ZN(new_n1132));
  AND4_X1   g706(.A1(new_n1131), .A2(new_n900), .A3(new_n901), .A4(new_n1132), .ZN(G308));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n900), .A3(new_n901), .A4(new_n1132), .ZN(G225));
endmodule


