

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590;

  XNOR2_X2 U321 ( .A(KEYINPUT48), .B(n412), .ZN(n452) );
  XNOR2_X1 U322 ( .A(n404), .B(n403), .ZN(n551) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n403) );
  NOR2_X1 U324 ( .A1(n531), .A2(n447), .ZN(n539) );
  XNOR2_X1 U325 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U326 ( .A(n381), .B(n363), .ZN(n366) );
  OR2_X1 U327 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U328 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U329 ( .A(n376), .B(n375), .ZN(n402) );
  INV_X1 U330 ( .A(G127GAT), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n461), .B(KEYINPUT120), .ZN(n462) );
  XNOR2_X1 U332 ( .A(n449), .B(KEYINPUT50), .ZN(n450) );
  XNOR2_X1 U333 ( .A(n463), .B(n462), .ZN(G1350GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U335 ( .A(G15GAT), .B(G1GAT), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n289), .B(KEYINPUT69), .ZN(n354) );
  XOR2_X1 U337 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n291) );
  XNOR2_X1 U338 ( .A(G8GAT), .B(G64GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n354), .B(n292), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n300) );
  XOR2_X1 U342 ( .A(G57GAT), .B(KEYINPUT72), .Z(n296) );
  XNOR2_X1 U343 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n394) );
  XOR2_X1 U345 ( .A(n394), .B(G155GAT), .Z(n298) );
  NAND2_X1 U346 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U349 ( .A(G211GAT), .B(G183GAT), .Z(n302) );
  XNOR2_X1 U350 ( .A(G22GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U352 ( .A(G78GAT), .B(n303), .ZN(n304) );
  XOR2_X1 U353 ( .A(n305), .B(n304), .Z(n466) );
  XOR2_X1 U354 ( .A(n466), .B(KEYINPUT105), .Z(n459) );
  XOR2_X1 U355 ( .A(G211GAT), .B(KEYINPUT21), .Z(n307) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n419) );
  XOR2_X1 U358 ( .A(G218GAT), .B(G162GAT), .Z(n372) );
  XOR2_X1 U359 ( .A(n419), .B(n372), .Z(n309) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U362 ( .A(n310), .B(G106GAT), .Z(n312) );
  XOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .Z(n356) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(n356), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT24), .B(KEYINPUT85), .Z(n314) );
  XNOR2_X1 U367 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT74), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n395) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n319), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X1 U375 ( .A(n395), .B(n432), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n471) );
  XOR2_X1 U377 ( .A(n471), .B(KEYINPUT66), .Z(n322) );
  XNOR2_X1 U378 ( .A(KEYINPUT28), .B(n322), .ZN(n531) );
  XOR2_X1 U379 ( .A(G134GAT), .B(G99GAT), .Z(n324) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G15GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U382 ( .A(G71GAT), .B(n325), .Z(n327) );
  NAND2_X1 U383 ( .A1(G227GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U385 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n329) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(G176GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U388 ( .A(n331), .B(n330), .Z(n341) );
  XOR2_X1 U389 ( .A(KEYINPUT81), .B(G127GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(G113GAT), .B(n334), .Z(n442) );
  XOR2_X1 U393 ( .A(G183GAT), .B(KEYINPUT83), .Z(n336) );
  XNOR2_X1 U394 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n337), .B(KEYINPUT18), .Z(n339) );
  XNOR2_X1 U397 ( .A(KEYINPUT84), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n416) );
  XNOR2_X1 U399 ( .A(n442), .B(n416), .ZN(n340) );
  XOR2_X1 U400 ( .A(n341), .B(n340), .Z(n528) );
  INV_X1 U401 ( .A(n528), .ZN(n478) );
  XOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n343) );
  NAND2_X1 U403 ( .A1(G229GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U405 ( .A(n344), .B(KEYINPUT30), .Z(n353) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n345), .B(G29GAT), .ZN(n346) );
  XOR2_X1 U408 ( .A(n346), .B(KEYINPUT8), .Z(n348) );
  XNOR2_X1 U409 ( .A(G43GAT), .B(G50GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n374) );
  XOR2_X1 U411 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n350) );
  XNOR2_X1 U412 ( .A(G197GAT), .B(G113GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n374), .B(n351), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n355) );
  XOR2_X1 U416 ( .A(n355), .B(n354), .Z(n358) );
  XOR2_X1 U417 ( .A(G169GAT), .B(G8GAT), .Z(n415) );
  XNOR2_X1 U418 ( .A(n356), .B(n415), .ZN(n357) );
  XOR2_X1 U419 ( .A(n358), .B(n357), .Z(n510) );
  XNOR2_X1 U420 ( .A(KEYINPUT71), .B(n510), .ZN(n559) );
  XOR2_X1 U421 ( .A(G85GAT), .B(G92GAT), .Z(n360) );
  XNOR2_X1 U422 ( .A(G99GAT), .B(G106GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n381) );
  NAND2_X1 U424 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  INV_X1 U425 ( .A(KEYINPUT9), .ZN(n361) );
  XOR2_X1 U426 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n365) );
  XNOR2_X1 U427 ( .A(G190GAT), .B(KEYINPUT11), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n367) );
  NAND2_X1 U429 ( .A1(n366), .A2(n367), .ZN(n371) );
  INV_X1 U430 ( .A(n366), .ZN(n369) );
  INV_X1 U431 ( .A(n367), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n369), .A2(n368), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n376) );
  XOR2_X1 U434 ( .A(G134GAT), .B(KEYINPUT78), .Z(n428) );
  XOR2_X1 U435 ( .A(n372), .B(n428), .Z(n373) );
  XOR2_X1 U436 ( .A(KEYINPUT79), .B(n402), .Z(n567) );
  XNOR2_X1 U437 ( .A(n567), .B(KEYINPUT36), .ZN(n494) );
  INV_X1 U438 ( .A(n466), .ZN(n585) );
  NAND2_X1 U439 ( .A1(n494), .A2(n585), .ZN(n379) );
  XOR2_X1 U440 ( .A(KEYINPUT45), .B(KEYINPUT107), .Z(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT65), .B(n377), .Z(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n398) );
  INV_X1 U443 ( .A(KEYINPUT32), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n383) );
  NAND2_X1 U445 ( .A1(G230GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n385) );
  INV_X1 U447 ( .A(KEYINPUT76), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U449 ( .A(G176GAT), .B(G64GAT), .Z(n413) );
  XNOR2_X1 U450 ( .A(G120GAT), .B(n413), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U452 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U455 ( .A1(n391), .A2(n390), .ZN(n393) );
  NAND2_X1 U456 ( .A1(n393), .A2(n392), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n404) );
  INV_X1 U459 ( .A(n404), .ZN(n580) );
  NOR2_X1 U460 ( .A1(n398), .A2(n580), .ZN(n399) );
  XOR2_X1 U461 ( .A(KEYINPUT108), .B(n399), .Z(n400) );
  NOR2_X1 U462 ( .A1(n559), .A2(n400), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n401), .B(KEYINPUT109), .ZN(n411) );
  BUF_X1 U464 ( .A(n402), .Z(n557) );
  INV_X1 U465 ( .A(n510), .ZN(n574) );
  NAND2_X1 U466 ( .A1(n574), .A2(n551), .ZN(n406) );
  XNOR2_X1 U467 ( .A(KEYINPUT106), .B(KEYINPUT46), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n407), .A2(n459), .ZN(n408) );
  NOR2_X1 U470 ( .A1(n557), .A2(n408), .ZN(n409) );
  XNOR2_X1 U471 ( .A(KEYINPUT47), .B(n409), .ZN(n410) );
  NAND2_X1 U472 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(G218GAT), .B(G92GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n424) );
  XOR2_X1 U475 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n422) );
  XNOR2_X1 U479 ( .A(G36GAT), .B(G204GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n486) );
  XNOR2_X1 U482 ( .A(KEYINPUT27), .B(n486), .ZN(n469) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G148GAT), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U486 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(n431), .B(KEYINPUT1), .Z(n434) );
  XNOR2_X1 U490 ( .A(n432), .B(KEYINPUT89), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U492 ( .A(KEYINPUT6), .B(G57GAT), .Z(n436) );
  XNOR2_X1 U493 ( .A(G141GAT), .B(G1GAT), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U495 ( .A(n438), .B(n437), .Z(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n440) );
  XNOR2_X1 U497 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n444), .B(n443), .Z(n475) );
  INV_X1 U501 ( .A(n475), .ZN(n522) );
  NAND2_X1 U502 ( .A1(n469), .A2(n522), .ZN(n445) );
  XOR2_X1 U503 ( .A(KEYINPUT90), .B(n445), .Z(n477) );
  NAND2_X1 U504 ( .A1(n452), .A2(n477), .ZN(n544) );
  NOR2_X1 U505 ( .A1(n478), .A2(n544), .ZN(n446) );
  XOR2_X1 U506 ( .A(KEYINPUT110), .B(n446), .Z(n447) );
  INV_X1 U507 ( .A(n539), .ZN(n448) );
  NOR2_X1 U508 ( .A1(n459), .A2(n448), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(G1342GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n454) );
  NAND2_X1 U511 ( .A1(n452), .A2(n486), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X2 U513 ( .A1(n455), .A2(n522), .ZN(n573) );
  NAND2_X1 U514 ( .A1(n471), .A2(n573), .ZN(n457) );
  INV_X1 U515 ( .A(KEYINPUT55), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X2 U517 ( .A1(n478), .A2(n458), .ZN(n568) );
  INV_X1 U518 ( .A(n568), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n460), .A2(n459), .ZN(n463) );
  INV_X1 U520 ( .A(G183GAT), .ZN(n461) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT93), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT34), .B(n465), .Z(n485) );
  NAND2_X1 U524 ( .A1(n559), .A2(n404), .ZN(n499) );
  NOR2_X1 U525 ( .A1(n567), .A2(n466), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT16), .ZN(n483) );
  NOR2_X1 U527 ( .A1(n528), .A2(n471), .ZN(n468) );
  XOR2_X1 U528 ( .A(n468), .B(KEYINPUT26), .Z(n545) );
  INV_X1 U529 ( .A(n545), .ZN(n572) );
  NAND2_X1 U530 ( .A1(n469), .A2(n572), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n528), .A2(n486), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n472), .Z(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n531), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT91), .B(n480), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n495) );
  NAND2_X1 U540 ( .A1(n483), .A2(n495), .ZN(n511) );
  NOR2_X1 U541 ( .A1(n499), .A2(n511), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n492), .A2(n522), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  BUF_X1 U544 ( .A(n486), .Z(n525) );
  NAND2_X1 U545 ( .A1(n525), .A2(n492), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT94), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n492), .A2(n528), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U552 ( .A1(n531), .A2(n492), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n494), .A2(n495), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n585), .A2(n496), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT96), .B(KEYINPUT37), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n521) );
  NOR2_X1 U558 ( .A1(n521), .A2(n499), .ZN(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT38), .B(n500), .ZN(n508) );
  NAND2_X1 U560 ( .A1(n508), .A2(n522), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT97), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n508), .A2(n525), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(KEYINPUT98), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n528), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  XOR2_X1 U573 ( .A(KEYINPUT99), .B(n551), .Z(n562) );
  NAND2_X1 U574 ( .A1(n510), .A2(n562), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n520), .A2(n511), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n522), .A2(n517), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n525), .A2(n517), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT100), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n528), .A2(n517), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n531), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  XOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT101), .Z(n524) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n532), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n532), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT102), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  XOR2_X1 U593 ( .A(G99GAT), .B(KEYINPUT103), .Z(n530) );
  NAND2_X1 U594 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT104), .Z(n534) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n535), .Z(G1339GAT) );
  NAND2_X1 U600 ( .A1(n539), .A2(n559), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n562), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n567), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT111), .Z(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT113), .Z(n547) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n574), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(n550), .Z(n553) );
  NAND2_X1 U618 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n556), .A2(n585), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n568), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .Z(n564) );
  NAND2_X1 U629 ( .A1(n568), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n576) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n587) );
  NAND2_X1 U639 ( .A1(n587), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(n577), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U645 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT124), .Z(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n585), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n494), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

