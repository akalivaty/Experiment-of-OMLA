//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G58), .B2(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(KEYINPUT67), .A2(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(KEYINPUT67), .A2(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n207), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n229), .C1(new_n218), .C2(new_n212), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  INV_X1    g0036(.A(G20), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g0039(.A1(new_n231), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT66), .Z(new_n241));
  NOR2_X1   g0041(.A1(new_n227), .A2(new_n241), .ZN(G361));
  XOR2_X1   g0042(.A(G226), .B(G232), .Z(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n255), .B(new_n256), .Z(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT69), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT69), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI211_X1 g0063(.A(G1), .B(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G232), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G226), .B2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n267), .A2(new_n272), .B1(new_n270), .B2(new_n217), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n264), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n274), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n224), .B2(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n281));
  XNOR2_X1  g0081(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n236), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n236), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n270), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n215), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n237), .A2(new_n270), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n222), .A2(new_n237), .B1(new_n202), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n277), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT73), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT12), .B1(new_n299), .B2(new_n222), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n285), .A2(new_n296), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n295), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n280), .A2(new_n281), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n307), .A2(G190), .A3(new_n308), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n283), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n282), .A2(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(G179), .A3(new_n308), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n282), .A2(new_n314), .A3(G169), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n310), .B1(new_n316), .B2(new_n306), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n288), .B1(new_n277), .B2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n203), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n319), .B1(new_n320), .B2(new_n292), .C1(new_n290), .C2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n318), .A2(G50), .B1(new_n288), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n298), .A2(new_n202), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n327));
  INV_X1    g0127(.A(new_n272), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G222), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n274), .C1(G77), .C2(new_n328), .ZN(new_n333));
  INV_X1    g0133(.A(new_n264), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n279), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n327), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT10), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n336), .A2(G179), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n325), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT15), .B(G87), .Z(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n321), .B(KEYINPUT71), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n292), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n284), .A2(new_n236), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n215), .B2(new_n298), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n215), .B2(new_n305), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n272), .A2(new_n330), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G238), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n211), .B2(new_n328), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n272), .A2(new_n265), .A3(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n274), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n276), .A2(G244), .A3(new_n278), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n334), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(G200), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n339), .B2(new_n360), .ZN(new_n362));
  AND4_X1   g0162(.A1(new_n317), .A2(new_n342), .A3(new_n346), .A4(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT74), .B1(new_n268), .B2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n270), .A3(KEYINPUT3), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n335), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(G223), .C2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n276), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n279), .A2(new_n265), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n372), .A2(new_n264), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G179), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n344), .B2(new_n374), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT78), .B1(new_n268), .B2(G33), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n270), .A3(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n380), .A3(new_n269), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n237), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT7), .A2(G20), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n272), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n383), .A2(new_n222), .A3(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(KEYINPUT67), .A2(G68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(KEYINPUT67), .A2(G68), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G58), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n237), .B1(new_n390), .B2(new_n233), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n292), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT76), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n201), .B1(new_n222), .B2(G58), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n237), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n377), .B1(new_n387), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n351), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT75), .B(new_n364), .C1(new_n365), .C2(new_n367), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n365), .A2(new_n367), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n269), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n384), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n366), .B1(KEYINPUT3), .B2(new_n270), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n268), .A2(KEYINPUT74), .A3(G33), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n269), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n410), .B2(new_n237), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(new_n412), .A3(G68), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n394), .A2(new_n398), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT77), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT77), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(new_n414), .A3(new_n417), .A4(KEYINPUT16), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n299), .A2(new_n321), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n318), .B2(new_n321), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n376), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT18), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(new_n418), .ZN(new_n425));
  INV_X1    g0225(.A(new_n401), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n374), .A2(G200), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n372), .A2(G190), .A3(new_n264), .A4(new_n373), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n435));
  NOR3_X1   g0235(.A1(new_n419), .A2(new_n432), .A3(new_n422), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n360), .A2(new_n344), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n353), .C1(G179), .C2(new_n360), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n363), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n404), .A2(G244), .A3(new_n330), .A4(new_n269), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n354), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n328), .A2(KEYINPUT4), .A3(G244), .A4(new_n330), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n274), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n260), .A2(new_n450), .A3(new_n261), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n263), .A2(G1), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n450), .A2(G41), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(G274), .A3(new_n276), .A4(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(KEYINPUT69), .A2(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT69), .A2(G41), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT5), .ZN(new_n461));
  INV_X1    g0261(.A(new_n453), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT81), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G257), .A3(new_n276), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n449), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G200), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n449), .A2(new_n339), .A3(new_n458), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n299), .A2(G97), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n383), .A2(G107), .A3(new_n386), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n292), .A2(new_n215), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n217), .A2(new_n211), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n237), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n472), .B1(new_n483), .B2(new_n351), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n286), .A2(new_n287), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n298), .B1(new_n277), .B2(G33), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n485), .B1(new_n484), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n471), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n467), .A2(G169), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n449), .A2(G179), .A3(new_n458), .A4(new_n466), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n472), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n385), .B1(new_n382), .B2(KEYINPUT7), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n474), .B(new_n481), .C1(new_n497), .C2(G107), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n489), .C1(new_n498), .C2(new_n285), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n224), .A2(new_n330), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n216), .A2(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n404), .A2(new_n269), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n276), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n462), .A2(new_n259), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n276), .A2(G250), .A3(new_n462), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G169), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n404), .A2(new_n237), .A3(G68), .A4(new_n269), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n289), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  NAND3_X1  g0313(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n237), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n478), .A2(new_n209), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n512), .A2(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n285), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n299), .A2(new_n347), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT82), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n488), .A2(new_n347), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n510), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G179), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n509), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n521), .A2(new_n523), .B1(G87), .B2(new_n488), .ZN(new_n529));
  NOR4_X1   g0329(.A1(new_n505), .A2(new_n508), .A3(new_n339), .A4(new_n506), .ZN(new_n530));
  INV_X1    g0330(.A(new_n509), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G200), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n526), .A2(new_n528), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n492), .A2(new_n500), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n465), .A2(G264), .A3(new_n276), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT90), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT90), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n465), .A2(new_n537), .A3(G264), .A4(new_n276), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n218), .A2(G1698), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n368), .B(new_n540), .C1(G250), .C2(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n276), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n539), .A2(new_n339), .A3(new_n458), .A4(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n463), .A2(G274), .A3(new_n457), .A4(new_n464), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n274), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n547), .B(new_n543), .C1(new_n536), .C2(new_n538), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n545), .B(KEYINPUT91), .C1(new_n548), .C2(G200), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT88), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n211), .B2(G20), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n211), .A2(KEYINPUT88), .A3(KEYINPUT23), .A4(G20), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n554), .B1(G116), .B2(new_n289), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n404), .A2(new_n237), .A3(G87), .A4(new_n269), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n237), .A3(G87), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT86), .A3(new_n269), .A4(new_n271), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT86), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n272), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n557), .A2(KEYINPUT87), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT87), .B1(new_n557), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n555), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(KEYINPUT24), .B(new_n555), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n351), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n488), .A2(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n299), .A2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(KEYINPUT25), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n576));
  MUX2_X1   g0376(.A(new_n573), .B(new_n575), .S(new_n576), .Z(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n548), .A2(KEYINPUT91), .A3(G200), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n534), .B1(new_n549), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n543), .B1(new_n536), .B2(new_n538), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n458), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n344), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n548), .A2(new_n527), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n487), .A2(G116), .A3(new_n285), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G283), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n237), .C1(G33), .C2(new_n217), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n351), .C1(new_n237), .C2(G116), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT20), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n587), .B1(G116), .B2(new_n299), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n465), .A2(G270), .A3(new_n276), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n218), .A2(new_n330), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n212), .A2(G1698), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n368), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n328), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n274), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n458), .A2(new_n596), .A3(new_n602), .A4(G190), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n458), .A2(new_n602), .A3(new_n596), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n595), .B(new_n603), .C1(new_n604), .C2(new_n468), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT85), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n458), .A2(new_n596), .A3(new_n602), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n594), .B1(new_n607), .B2(G200), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n603), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n458), .A2(new_n596), .A3(new_n602), .A4(G179), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n595), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT84), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n607), .A2(G169), .A3(new_n594), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n611), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n581), .A2(new_n586), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n442), .A2(new_n623), .ZN(G372));
  NAND3_X1  g0424(.A1(new_n586), .A2(new_n615), .A3(new_n620), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n492), .A2(new_n500), .A3(new_n533), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n571), .A2(new_n572), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n583), .A2(new_n628), .A3(new_n468), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(new_n577), .A3(new_n549), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n523), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n525), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n634), .B(new_n528), .C1(G169), .C2(new_n509), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n495), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n495), .A2(new_n636), .A3(KEYINPUT92), .A4(new_n637), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n533), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n532), .A2(new_n529), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT26), .B1(new_n645), .B2(new_n500), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n631), .A2(new_n635), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n441), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n346), .ZN(new_n649));
  INV_X1    g0449(.A(new_n437), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n316), .A2(new_n306), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n310), .A2(new_n440), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n423), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(new_n342), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(G369));
  NAND2_X1  g0459(.A1(new_n615), .A2(new_n620), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n297), .A2(G20), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n277), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(KEYINPUT93), .B(G343), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n578), .A2(new_n668), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT94), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT94), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n578), .A2(new_n674), .A3(new_n668), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n630), .A3(new_n586), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT95), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT95), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n580), .A2(new_n549), .B1(new_n672), .B2(KEYINPUT94), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n586), .A2(new_n675), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n671), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT96), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n586), .A2(new_n668), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n676), .A2(KEYINPUT95), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n679), .A2(new_n680), .A3(new_n678), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n670), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT96), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n668), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n687), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n595), .A2(new_n669), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n660), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n621), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n691), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n262), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n229), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n516), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n235), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n647), .A2(new_n669), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n494), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n582), .A3(new_n509), .A4(new_n604), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n539), .A2(new_n544), .A3(new_n509), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n714), .A4(new_n604), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n607), .A2(new_n527), .A3(new_n531), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT97), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n607), .A2(new_n531), .A3(KEYINPUT97), .A4(new_n527), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n583), .A3(new_n467), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n668), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n623), .B2(new_n668), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(new_n635), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n645), .A2(new_n500), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n641), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n640), .A2(new_n533), .A3(new_n642), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n631), .B(new_n733), .C1(new_n641), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n669), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n713), .A2(new_n730), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n710), .B1(new_n738), .B2(G1), .ZN(G364));
  INV_X1    g0539(.A(new_n699), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n277), .B1(new_n661), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n704), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n698), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n236), .B1(G20), .B2(new_n344), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n468), .A2(G179), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G20), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n237), .B1(new_n752), .B2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(G303), .B1(new_n754), .B2(G294), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n237), .A2(new_n527), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G326), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n272), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n750), .A2(new_n527), .A3(G200), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n761), .A2(G322), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n237), .A2(G190), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(new_n752), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(G329), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n756), .A2(new_n339), .A3(G200), .ZN(new_n766));
  OR2_X1    g0566(.A1(KEYINPUT33), .A2(G317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(KEYINPUT33), .A2(G317), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n760), .A2(new_n762), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n527), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G311), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n748), .A2(new_n763), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n770), .B(new_n774), .C1(new_n775), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT99), .ZN(new_n781));
  INV_X1    g0581(.A(new_n764), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT32), .B1(new_n782), .B2(new_n392), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n202), .B2(new_n757), .ZN(new_n784));
  INV_X1    g0584(.A(new_n761), .ZN(new_n785));
  INV_X1    g0585(.A(G58), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n786), .B1(new_n772), .B2(new_n215), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n782), .A2(KEYINPUT32), .A3(new_n392), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n766), .A2(new_n304), .B1(new_n753), .B2(new_n217), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G87), .B2(new_n751), .ZN(new_n791));
  INV_X1    g0591(.A(new_n779), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G107), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n789), .A2(new_n328), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n747), .B1(new_n781), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n746), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n229), .A2(new_n272), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G355), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n410), .A2(KEYINPUT75), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n368), .A2(new_n403), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n229), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G45), .B2(new_n708), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n254), .A2(G45), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n801), .B1(G116), .B2(new_n228), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n795), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n798), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n743), .B(new_n810), .C1(new_n698), .C2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n745), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n353), .A2(new_n668), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n362), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n440), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n440), .A2(new_n668), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n692), .A2(new_n660), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n493), .A2(new_n494), .B1(new_n484), .B2(new_n489), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n636), .A2(new_n637), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n471), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n629), .A2(new_n572), .A3(new_n571), .A4(new_n577), .ZN(new_n826));
  INV_X1    g0626(.A(new_n549), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n533), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n646), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n643), .A2(new_n635), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n669), .B(new_n821), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n647), .A2(KEYINPUT101), .A3(new_n669), .A4(new_n821), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(new_n711), .B2(new_n820), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(new_n730), .Z(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n743), .ZN(new_n837));
  INV_X1    g0637(.A(new_n743), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n820), .B2(new_n796), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n757), .A2(new_n600), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n785), .A2(new_n841), .B1(new_n766), .B2(new_n775), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G107), .C2(new_n751), .ZN(new_n843));
  INV_X1    g0643(.A(G116), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n772), .A2(new_n844), .B1(new_n753), .B2(new_n217), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n328), .B(new_n845), .C1(G311), .C2(new_n764), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(new_n209), .C2(new_n779), .ZN(new_n847));
  INV_X1    g0647(.A(new_n766), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n758), .B1(new_n848), .B2(G150), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n761), .A2(G143), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(new_n392), .C2(new_n772), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n851), .A2(new_n852), .B1(G50), .B2(new_n751), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n792), .A2(G68), .B1(G132), .B2(new_n764), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n853), .A2(new_n854), .A3(new_n805), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n753), .A2(new_n786), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n746), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n746), .A2(new_n796), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n839), .B(new_n859), .C1(G77), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT100), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n837), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  INV_X1    g0665(.A(KEYINPUT105), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n413), .A2(new_n414), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n486), .B1(new_n868), .B2(new_n377), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n411), .B1(new_n804), .B2(new_n384), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n399), .B1(new_n870), .B2(G68), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n417), .B1(new_n871), .B2(KEYINPUT16), .ZN(new_n872));
  INV_X1    g0672(.A(new_n418), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n421), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(new_n376), .B1(new_n427), .B2(new_n433), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n665), .B1(new_n874), .B2(new_n421), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n867), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n436), .ZN(new_n880));
  INV_X1    g0680(.A(new_n665), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n419), .A2(new_n422), .B1(new_n376), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n866), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n877), .B1(new_n424), .B2(new_n437), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(new_n376), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n874), .B2(new_n421), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n877), .A2(new_n889), .A3(new_n436), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT105), .B(new_n887), .C1(new_n890), .C2(new_n867), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n885), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n891), .A4(new_n886), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR4_X1   g0696(.A1(new_n828), .A2(new_n692), .A3(new_n621), .A4(new_n668), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n725), .A2(new_n668), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT31), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT107), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT107), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n728), .B(new_n904), .C1(new_n623), .C2(new_n668), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n820), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n306), .A2(new_n668), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n652), .A2(new_n668), .B1(new_n317), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n896), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n820), .B(new_n908), .C1(new_n903), .C2(new_n905), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT108), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n881), .B1(new_n419), .B2(new_n422), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n650), .B2(new_n656), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n883), .B1(new_n880), .B2(new_n882), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n884), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n893), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n914), .B1(new_n895), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n895), .A2(new_n914), .A3(new_n919), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n913), .B(KEYINPUT40), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n912), .A2(new_n922), .A3(G330), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n903), .A2(new_n905), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n441), .A2(G330), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n895), .A2(new_n919), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT108), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n895), .A2(new_n914), .A3(new_n919), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n911), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n913), .B1(new_n910), .B2(new_n911), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n441), .A3(new_n924), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n646), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n581), .B2(new_n625), .ZN(new_n936));
  INV_X1    g0736(.A(new_n830), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n668), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT101), .B1(new_n938), .B2(new_n821), .ZN(new_n939));
  INV_X1    g0739(.A(new_n834), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n819), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT103), .A3(new_n909), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT103), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n818), .B1(new_n833), .B2(new_n834), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n908), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n945), .A3(new_n896), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n894), .B2(new_n895), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n895), .A2(new_n947), .A3(new_n919), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n651), .A2(KEYINPUT106), .A3(new_n668), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT106), .B1(new_n651), .B2(new_n668), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n424), .A2(new_n665), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n946), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n737), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n441), .B1(new_n957), .B2(new_n712), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n658), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n956), .B(new_n959), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n934), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n277), .B2(new_n661), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n479), .A2(new_n480), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT102), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n844), .B1(new_n964), .B2(KEYINPUT35), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n965), .B(new_n238), .C1(KEYINPUT35), .C2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n235), .A2(G77), .A3(new_n390), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(G50), .B2(new_n304), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n297), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n967), .A3(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n825), .B1(new_n824), .B2(new_n669), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n638), .A2(new_n669), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT42), .B1(new_n682), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n977), .C1(new_n689), .C2(new_n684), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n823), .A2(new_n669), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n529), .A2(new_n669), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT110), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n731), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT111), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n645), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n983), .B2(new_n985), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n976), .A2(new_n978), .A3(new_n991), .A4(new_n979), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n983), .A2(KEYINPUT43), .A3(new_n985), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n990), .A2(KEYINPUT112), .A3(new_n992), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n701), .A2(new_n975), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n704), .B(KEYINPUT41), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n975), .B1(new_n686), .B2(new_n690), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n686), .A2(new_n690), .A3(new_n975), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT44), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n700), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1003), .B(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1006), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n701), .A3(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n682), .A2(KEYINPUT113), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n682), .B(KEYINPUT113), .C1(new_n694), .C2(new_n671), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n740), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n699), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n738), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1008), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n738), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n741), .B(KEYINPUT114), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n1000), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n758), .A2(G311), .B1(new_n754), .B2(G107), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n751), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n844), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1026), .A2(KEYINPUT46), .B1(G303), .B2(new_n761), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(KEYINPUT46), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1024), .B(new_n1027), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n805), .B1(G294), .B2(new_n848), .ZN(new_n1033));
  INV_X1    g0833(.A(G317), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n775), .B2(new_n772), .C1(new_n1034), .C2(new_n782), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n776), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1032), .B(new_n1035), .C1(G97), .C2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G143), .A2(new_n758), .B1(new_n848), .B2(G159), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n202), .B2(new_n772), .C1(new_n786), .C2(new_n1025), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT116), .B(G137), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n764), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n215), .B2(new_n776), .C1(new_n320), .C2(new_n785), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G68), .B2(new_n754), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1037), .B1(new_n1043), .B2(new_n328), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT47), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n746), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n983), .A2(new_n985), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n798), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n347), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n806), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n799), .B1(new_n228), .B2(new_n1049), .C1(new_n1050), .C2(new_n250), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n743), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1023), .A2(new_n1052), .ZN(G387));
  NAND3_X1  g0853(.A1(new_n1016), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n247), .A2(new_n263), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n706), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1055), .A2(new_n806), .B1(new_n1056), .B2(new_n800), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n349), .A2(G50), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT50), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n263), .B1(new_n304), .B2(new_n215), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1059), .A2(new_n1056), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1057), .A2(new_n1061), .B1(G107), .B2(new_n228), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n838), .B1(new_n1062), .B2(new_n799), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT117), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n848), .B1(new_n758), .B2(G322), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n600), .B2(new_n772), .C1(new_n1034), .C2(new_n785), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT48), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n775), .B2(new_n753), .C1(new_n841), .C2(new_n1025), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n805), .B1(G326), .B2(new_n764), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n844), .C2(new_n776), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1025), .A2(new_n215), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n792), .A2(G97), .B1(G150), .B2(new_n764), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n304), .B2(new_n772), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G50), .C2(new_n761), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n321), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n848), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n758), .A2(G159), .B1(new_n754), .B2(new_n347), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n805), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1064), .B1(new_n694), .B2(new_n811), .C1(new_n1081), .C2(new_n747), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n738), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(new_n705), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1054), .B(new_n1082), .C1(new_n1084), .C2(new_n1019), .ZN(G393));
  NAND3_X1  g0885(.A1(new_n1008), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n838), .B1(new_n975), .B2(new_n798), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n799), .B1(new_n217), .B2(new_n228), .C1(new_n1050), .C2(new_n257), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n758), .A2(G317), .B1(G311), .B2(new_n761), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G294), .B2(new_n773), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n764), .A2(G322), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1025), .A2(new_n775), .B1(new_n753), .B2(new_n844), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G303), .B2(new_n848), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n328), .B1(new_n792), .B2(G107), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n758), .A2(G150), .B1(G159), .B2(new_n761), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G87), .B2(new_n792), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n349), .A2(new_n772), .B1(new_n202), .B2(new_n766), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n753), .A2(new_n215), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n804), .B1(G143), .B2(new_n764), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1025), .A2(new_n223), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1096), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n746), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1087), .A2(new_n1088), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n705), .B1(new_n1110), .B2(new_n1018), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1111), .B2(new_n1020), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  NAND3_X1  g0913(.A1(new_n958), .A2(new_n925), .A3(new_n658), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n908), .B1(new_n730), .B2(new_n820), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n906), .A2(new_n909), .ZN(new_n1116));
  INV_X1    g0916(.A(G330), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n941), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n735), .A2(new_n669), .A3(new_n817), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n819), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n730), .A2(new_n820), .A3(new_n908), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n906), .A2(G330), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1122), .B(new_n1124), .C1(new_n1125), .C2(new_n909), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1114), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n953), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n944), .B2(new_n908), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n948), .A2(new_n949), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1121), .A2(new_n909), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n953), .B(KEYINPUT119), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n921), .C2(new_n920), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1131), .A2(new_n1123), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1127), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT120), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1114), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(KEYINPUT120), .B(new_n1114), .C1(new_n1119), .C2(new_n1126), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n704), .B(new_n1138), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n950), .A2(new_n797), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n751), .A2(G87), .B1(new_n764), .B2(G294), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n211), .B2(new_n766), .C1(new_n775), .C2(new_n757), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1101), .B(new_n1149), .C1(G97), .C2(new_n773), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n844), .B2(new_n785), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n328), .B(new_n1151), .C1(G68), .C2(new_n792), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT121), .Z(new_n1153));
  AOI22_X1  g0953(.A1(new_n758), .A2(G128), .B1(new_n754), .B2(G159), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n848), .A2(new_n1040), .ZN(new_n1155));
  INV_X1    g0955(.A(G132), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1155), .C1(new_n1156), .C2(new_n785), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT54), .B(G143), .Z(new_n1158));
  AOI211_X1 g0958(.A(new_n272), .B(new_n1157), .C1(new_n773), .C2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n764), .A2(G125), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n202), .C2(new_n776), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n751), .A2(G150), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT122), .Z(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(new_n747), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1147), .A2(new_n838), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1077), .B2(new_n861), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1022), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT123), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT123), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1146), .B1(new_n1170), .B2(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n342), .A2(new_n346), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n325), .A2(new_n881), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n796), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1036), .A2(G58), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n844), .B2(new_n757), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n804), .A2(new_n262), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G68), .C2(new_n754), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1049), .A2(new_n772), .B1(new_n785), .B2(new_n211), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1184), .B(new_n1073), .C1(G283), .C2(new_n764), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(new_n217), .C2(new_n766), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT58), .Z(new_n1187));
  OAI211_X1 g0987(.A(new_n1182), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n848), .A2(G132), .B1(new_n773), .B2(G137), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n751), .A2(new_n1158), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n758), .A2(G125), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n754), .A2(G150), .B1(G128), .B2(new_n761), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT59), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n392), .B2(new_n776), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1188), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n746), .B1(new_n1187), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n860), .A2(new_n202), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1179), .A2(new_n743), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n946), .A2(new_n954), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n932), .A2(G330), .A3(new_n1177), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n923), .A2(new_n1178), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n955), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1177), .B1(new_n932), .B2(G330), .ZN(new_n1206));
  AND4_X1   g1006(.A1(G330), .A2(new_n912), .A3(new_n922), .A4(new_n1177), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n956), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1201), .B1(new_n1209), .B2(new_n1022), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1205), .A2(new_n1208), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n704), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1212), .B2(new_n1216), .ZN(G375));
  NOR2_X1   g1017(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1144), .A2(new_n1002), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n772), .A2(new_n211), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1025), .A2(new_n217), .B1(new_n757), .B2(new_n841), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G116), .C2(new_n848), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n782), .A2(new_n600), .B1(new_n1049), .B2(new_n753), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n328), .B(new_n1223), .C1(G283), .C2(new_n761), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n215), .C2(new_n779), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n805), .B1(new_n1226), .B2(new_n782), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n772), .A2(new_n320), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n757), .A2(new_n1156), .B1(new_n753), .B2(new_n202), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G159), .C2(new_n751), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n848), .A2(new_n1158), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n761), .A2(new_n1040), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n1180), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n746), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n743), .B(new_n1235), .C1(new_n909), .C2(new_n797), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n304), .B2(new_n860), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1140), .B2(new_n1022), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1219), .A2(new_n1238), .ZN(G381));
  NAND3_X1  g1039(.A1(new_n1146), .A2(new_n1169), .A3(new_n1168), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G375), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G381), .A2(G384), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1023), .A2(new_n1052), .A3(new_n1112), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1241), .B2(new_n667), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G407), .ZN(G409));
  NOR2_X1   g1048(.A1(new_n666), .A2(new_n1246), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(G2897), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT126), .Z(new_n1251));
  NAND2_X1  g1051(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1127), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n704), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1238), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n705), .B1(new_n1218), .B2(KEYINPUT60), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1258), .B(new_n1253), .C1(KEYINPUT60), .C2(new_n1218), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1259), .B2(new_n1238), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1251), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1238), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n864), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1251), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1256), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1209), .A2(new_n1001), .A3(new_n1213), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1209), .A2(new_n1213), .A3(KEYINPUT124), .A4(new_n1001), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1210), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1240), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1210), .C1(new_n1212), .C2(new_n1216), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1249), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1266), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n813), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1112), .B1(new_n1023), .B2(new_n1052), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1243), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(G390), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1023), .A2(new_n1052), .A3(new_n1112), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1278), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1280), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1280), .A2(new_n1284), .A3(KEYINPUT127), .A4(new_n1285), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1277), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1263), .A2(new_n1256), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1249), .B(new_n1291), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1292), .B2(KEYINPUT63), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1291), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1275), .A2(new_n1276), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(KEYINPUT125), .A3(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1290), .A2(new_n1293), .A3(new_n1295), .A4(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1257), .A2(new_n1260), .A3(new_n1251), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1264), .B1(new_n1263), .B2(new_n1256), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1209), .A2(new_n1022), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1200), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n705), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1211), .A2(KEYINPUT57), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1309), .A2(G378), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1310), .B2(new_n1249), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT62), .B1(new_n1311), .B2(new_n1297), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1285), .B1(new_n1292), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1301), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1300), .A2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1272), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1301), .A2(new_n1274), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1274), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1291), .ZN(G402));
endmodule


