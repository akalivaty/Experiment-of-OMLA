

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n677), .A2(n676), .ZN(n727) );
  INV_X1 U551 ( .A(G2104), .ZN(n520) );
  AND2_X1 U552 ( .A1(G125), .A2(n872), .ZN(n513) );
  INV_X1 U553 ( .A(n727), .ZN(n679) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n684) );
  XNOR2_X1 U555 ( .A(n712), .B(KEYINPUT30), .ZN(n713) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n717) );
  AND2_X1 U557 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U558 ( .A1(G8), .A2(n727), .ZN(n756) );
  XNOR2_X1 U559 ( .A(n521), .B(KEYINPUT65), .ZN(n872) );
  NOR2_X1 U560 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U561 ( .A1(G651), .A2(n607), .ZN(n636) );
  AND2_X1 U562 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U563 ( .A(n525), .B(KEYINPUT64), .ZN(G160) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n514), .Z(n866) );
  NAND2_X1 U566 ( .A1(G137), .A2(n866), .ZN(n517) );
  NAND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XOR2_X2 U568 ( .A(KEYINPUT66), .B(n515), .Z(n870) );
  NAND2_X1 U569 ( .A1(G113), .A2(n870), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U571 ( .A(n518), .B(KEYINPUT67), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G2105), .A2(n520), .ZN(n867) );
  NAND2_X1 U573 ( .A1(G101), .A2(n867), .ZN(n519) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(n519), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n520), .A2(G2105), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n522), .A2(n513), .ZN(n523) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n629) );
  NAND2_X1 U578 ( .A1(G85), .A2(n629), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n607) );
  INV_X1 U580 ( .A(G651), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n607), .A2(n528), .ZN(n627) );
  NAND2_X1 U582 ( .A1(G72), .A2(n627), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n636), .A2(G47), .ZN(n533) );
  NOR2_X1 U585 ( .A1(G543), .A2(n528), .ZN(n530) );
  XNOR2_X1 U586 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n529) );
  XNOR2_X1 U587 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U588 ( .A(KEYINPUT68), .B(n531), .ZN(n633) );
  NAND2_X1 U589 ( .A1(G60), .A2(n633), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  OR2_X1 U591 ( .A1(n535), .A2(n534), .ZN(G290) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  NAND2_X1 U594 ( .A1(n636), .A2(G52), .ZN(n537) );
  NAND2_X1 U595 ( .A1(G64), .A2(n633), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U597 ( .A(KEYINPUT70), .B(n538), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G90), .A2(n629), .ZN(n540) );
  NAND2_X1 U599 ( .A1(G77), .A2(n627), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U601 ( .A(KEYINPUT9), .B(n541), .ZN(n542) );
  XNOR2_X1 U602 ( .A(KEYINPUT71), .B(n542), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n544), .A2(n543), .ZN(G171) );
  NAND2_X1 U604 ( .A1(n636), .A2(G51), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G63), .A2(n633), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U607 ( .A(KEYINPUT6), .B(n547), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n629), .A2(G89), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G76), .A2(n627), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U612 ( .A(n551), .B(KEYINPUT5), .Z(n552) );
  NOR2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT77), .B(n554), .Z(n555) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(n555), .Z(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n558) );
  INV_X1 U620 ( .A(G223), .ZN(n810) );
  NAND2_X1 U621 ( .A1(G567), .A2(n810), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(G234) );
  NAND2_X1 U623 ( .A1(n633), .A2(G56), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n559), .Z(n565) );
  NAND2_X1 U625 ( .A1(n629), .A2(G81), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G68), .A2(n627), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n636), .A2(G43), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n908) );
  INV_X1 U633 ( .A(n908), .ZN(n641) );
  NAND2_X1 U634 ( .A1(n641), .A2(G860), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n629), .A2(G92), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G66), .A2(n633), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n627), .A2(G79), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT75), .B(n570), .Z(n572) );
  NAND2_X1 U642 ( .A1(n636), .A2(G54), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U644 ( .A(KEYINPUT76), .B(n573), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT15), .ZN(n917) );
  INV_X1 U647 ( .A(G868), .ZN(n650) );
  NAND2_X1 U648 ( .A1(n917), .A2(n650), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U650 ( .A1(n636), .A2(G53), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G65), .A2(n633), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G91), .A2(n629), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G78), .A2(n627), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n907) );
  INV_X1 U657 ( .A(n907), .ZN(G299) );
  XNOR2_X1 U658 ( .A(KEYINPUT78), .B(n650), .ZN(n585) );
  NOR2_X1 U659 ( .A1(G286), .A2(n585), .ZN(n587) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(G297) );
  INV_X1 U662 ( .A(G860), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n588), .A2(G559), .ZN(n589) );
  INV_X1 U664 ( .A(n917), .ZN(n648) );
  NAND2_X1 U665 ( .A1(n589), .A2(n648), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G868), .A2(n908), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G868), .A2(n648), .ZN(n591) );
  NOR2_X1 U669 ( .A1(G559), .A2(n591), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U671 ( .A(KEYINPUT79), .B(n594), .Z(G282) );
  NAND2_X1 U672 ( .A1(G135), .A2(n866), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n595), .B(KEYINPUT80), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G123), .A2(n872), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U676 ( .A1(G111), .A2(n870), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U678 ( .A1(G99), .A2(n867), .ZN(n599) );
  XNOR2_X1 U679 ( .A(KEYINPUT81), .B(n599), .ZN(n600) );
  NOR2_X1 U680 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n936) );
  XNOR2_X1 U682 ( .A(G2096), .B(n936), .ZN(n604) );
  NOR2_X1 U683 ( .A1(G2100), .A2(n604), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT82), .B(n605), .Z(G156) );
  NAND2_X1 U685 ( .A1(G49), .A2(n636), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT88), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G87), .A2(n607), .ZN(n608) );
  XOR2_X1 U688 ( .A(KEYINPUT89), .B(n608), .Z(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n633), .A2(n611), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G651), .A2(G74), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G288) );
  NAND2_X1 U693 ( .A1(G88), .A2(n629), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G75), .A2(n627), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n636), .A2(G50), .ZN(n617) );
  NAND2_X1 U697 ( .A1(G62), .A2(n633), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U699 ( .A1(n619), .A2(n618), .ZN(G166) );
  NAND2_X1 U700 ( .A1(n629), .A2(G86), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G61), .A2(n633), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n627), .A2(G73), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n636), .A2(G48), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U708 ( .A1(n627), .A2(G80), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(KEYINPUT84), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G93), .A2(n629), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(KEYINPUT85), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G67), .A2(n633), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n636), .A2(G55), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT86), .B(n637), .Z(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U718 ( .A(KEYINPUT87), .B(n640), .ZN(n822) );
  XNOR2_X1 U719 ( .A(n822), .B(n641), .ZN(n647) );
  XNOR2_X1 U720 ( .A(G166), .B(KEYINPUT19), .ZN(n643) );
  XNOR2_X1 U721 ( .A(G290), .B(n907), .ZN(n642) );
  XNOR2_X1 U722 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U723 ( .A(n644), .B(G305), .Z(n645) );
  XNOR2_X1 U724 ( .A(G288), .B(n645), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n647), .B(n646), .ZN(n884) );
  NAND2_X1 U726 ( .A1(n648), .A2(G559), .ZN(n818) );
  XOR2_X1 U727 ( .A(n884), .B(n818), .Z(n649) );
  NAND2_X1 U728 ( .A1(G868), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n822), .A2(n650), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n653) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n653), .Z(n654) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(n655), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n656), .A2(G2072), .ZN(G158) );
  XOR2_X1 U736 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U738 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NAND2_X1 U739 ( .A1(G69), .A2(G120), .ZN(n657) );
  NOR2_X1 U740 ( .A1(G237), .A2(n657), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G108), .A2(n658), .ZN(n816) );
  NAND2_X1 U742 ( .A1(G567), .A2(n816), .ZN(n663) );
  NOR2_X1 U743 ( .A1(G219), .A2(G220), .ZN(n659) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U745 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(G96), .A2(n661), .ZN(n817) );
  NAND2_X1 U747 ( .A1(G2106), .A2(n817), .ZN(n662) );
  NAND2_X1 U748 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U749 ( .A(KEYINPUT90), .B(n664), .Z(G319) );
  INV_X1 U750 ( .A(G319), .ZN(n666) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n665) );
  NOR2_X1 U752 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U753 ( .A(KEYINPUT91), .B(n667), .Z(n815) );
  NAND2_X1 U754 ( .A1(n815), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(G138), .A2(n866), .ZN(n669) );
  NAND2_X1 U756 ( .A1(G102), .A2(n867), .ZN(n668) );
  NAND2_X1 U757 ( .A1(n669), .A2(n668), .ZN(n674) );
  NAND2_X1 U758 ( .A1(G126), .A2(n872), .ZN(n670) );
  XNOR2_X1 U759 ( .A(n670), .B(KEYINPUT92), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G114), .A2(n870), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U762 ( .A1(n674), .A2(n673), .ZN(G164) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U764 ( .A(G1986), .B(G290), .ZN(n914) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G40), .A2(G160), .ZN(n675) );
  NOR2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n804) );
  NAND2_X1 U768 ( .A1(n914), .A2(n804), .ZN(n792) );
  INV_X1 U769 ( .A(n675), .ZN(n677) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n756), .ZN(n722) );
  INV_X1 U771 ( .A(n727), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G1956), .B(KEYINPUT97), .ZN(n986) );
  NOR2_X1 U773 ( .A1(n705), .A2(n986), .ZN(n678) );
  XNOR2_X1 U774 ( .A(KEYINPUT98), .B(n678), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n679), .A2(G2072), .ZN(n680) );
  XNOR2_X1 U776 ( .A(n680), .B(KEYINPUT27), .ZN(n681) );
  XNOR2_X1 U777 ( .A(n681), .B(KEYINPUT96), .ZN(n682) );
  NOR2_X1 U778 ( .A1(n683), .A2(n682), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n907), .A2(n686), .ZN(n685) );
  XNOR2_X1 U780 ( .A(n685), .B(n684), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n907), .A2(n686), .ZN(n699) );
  INV_X1 U782 ( .A(G1996), .ZN(n960) );
  NOR2_X1 U783 ( .A1(n727), .A2(n960), .ZN(n687) );
  XOR2_X1 U784 ( .A(n687), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U785 ( .A1(n727), .A2(G1341), .ZN(n688) );
  NAND2_X1 U786 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U787 ( .A1(n908), .A2(n690), .ZN(n694) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n727), .ZN(n692) );
  NAND2_X1 U789 ( .A1(G2067), .A2(n705), .ZN(n691) );
  NAND2_X1 U790 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n917), .A2(n695), .ZN(n693) );
  OR2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n917), .A2(n695), .ZN(n696) );
  NAND2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U797 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n703), .B(n702), .ZN(n709) );
  OR2_X1 U799 ( .A1(n705), .A2(G1961), .ZN(n707) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT95), .Z(n704) );
  XNOR2_X1 U801 ( .A(KEYINPUT25), .B(n704), .ZN(n959) );
  NAND2_X1 U802 ( .A1(n705), .A2(n959), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n714), .A2(G171), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n720) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n727), .ZN(n723) );
  NOR2_X1 U807 ( .A1(n722), .A2(n723), .ZN(n710) );
  XNOR2_X1 U808 ( .A(KEYINPUT100), .B(n710), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n711), .A2(G8), .ZN(n712) );
  NOR2_X1 U810 ( .A1(n713), .A2(G168), .ZN(n716) );
  NOR2_X1 U811 ( .A1(G171), .A2(n714), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U813 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n726) );
  INV_X1 U815 ( .A(n726), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U817 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n738) );
  NAND2_X1 U819 ( .A1(n726), .A2(G286), .ZN(n734) );
  INV_X1 U820 ( .A(G8), .ZN(n732) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n756), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U826 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n735) );
  XNOR2_X1 U827 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n752) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n924) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n739) );
  XNOR2_X1 U831 ( .A(KEYINPUT102), .B(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n924), .A2(n740), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n752), .A2(n741), .ZN(n744) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n921) );
  INV_X1 U835 ( .A(n921), .ZN(n742) );
  NOR2_X1 U836 ( .A1(n756), .A2(n742), .ZN(n743) );
  AND2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U838 ( .A1(KEYINPUT33), .A2(n745), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n924), .A2(KEYINPUT33), .ZN(n746) );
  NOR2_X1 U840 ( .A1(n746), .A2(n756), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n904) );
  NAND2_X1 U843 ( .A1(n749), .A2(n904), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U845 ( .A1(G8), .A2(n750), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U847 ( .A1(n753), .A2(n756), .ZN(n758) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n754) );
  XOR2_X1 U849 ( .A(n754), .B(KEYINPUT24), .Z(n755) );
  NOR2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n790) );
  NAND2_X1 U853 ( .A1(G131), .A2(n866), .ZN(n762) );
  NAND2_X1 U854 ( .A1(G95), .A2(n867), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n872), .A2(G119), .ZN(n763) );
  XOR2_X1 U857 ( .A(KEYINPUT94), .B(n763), .Z(n764) );
  NOR2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n767) );
  NAND2_X1 U859 ( .A1(G107), .A2(n870), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n862) );
  AND2_X1 U861 ( .A1(n862), .A2(G1991), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G141), .A2(n866), .ZN(n769) );
  NAND2_X1 U863 ( .A1(G129), .A2(n872), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n867), .A2(G105), .ZN(n770) );
  XOR2_X1 U866 ( .A(KEYINPUT38), .B(n770), .Z(n771) );
  NOR2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U868 ( .A1(G117), .A2(n870), .ZN(n773) );
  NAND2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n859) );
  AND2_X1 U870 ( .A1(n859), .A2(G1996), .ZN(n775) );
  NOR2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n937) );
  INV_X1 U872 ( .A(n804), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n937), .A2(n777), .ZN(n795) );
  INV_X1 U874 ( .A(n795), .ZN(n788) );
  XNOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NAND2_X1 U876 ( .A1(n872), .A2(G128), .ZN(n778) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(n778), .Z(n780) );
  NAND2_X1 U878 ( .A1(G116), .A2(n870), .ZN(n779) );
  NAND2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U880 ( .A(n781), .B(KEYINPUT35), .ZN(n786) );
  NAND2_X1 U881 ( .A1(G140), .A2(n866), .ZN(n783) );
  NAND2_X1 U882 ( .A1(G104), .A2(n867), .ZN(n782) );
  NAND2_X1 U883 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U884 ( .A(KEYINPUT34), .B(n784), .Z(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U886 ( .A(n787), .B(KEYINPUT36), .Z(n881) );
  NOR2_X1 U887 ( .A1(n801), .A2(n881), .ZN(n947) );
  NAND2_X1 U888 ( .A1(n804), .A2(n947), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n788), .A2(n799), .ZN(n789) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n807) );
  XOR2_X1 U891 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n798) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n859), .ZN(n941) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n793) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n862), .ZN(n939) );
  NOR2_X1 U895 ( .A1(n793), .A2(n939), .ZN(n794) );
  NOR2_X1 U896 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U897 ( .A1(n941), .A2(n796), .ZN(n797) );
  XNOR2_X1 U898 ( .A(n798), .B(n797), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n803) );
  AND2_X1 U900 ( .A1(n801), .A2(n881), .ZN(n802) );
  XOR2_X1 U901 ( .A(KEYINPUT104), .B(n802), .Z(n951) );
  NAND2_X1 U902 ( .A1(n803), .A2(n951), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n808) );
  XNOR2_X1 U906 ( .A(n809), .B(n808), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n810), .ZN(G217) );
  NAND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n812) );
  INV_X1 U909 ( .A(G661), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U911 ( .A(n813), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(G188) );
  XOR2_X1 U914 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  XNOR2_X1 U915 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(G325) );
  XOR2_X1 U917 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U919 ( .A(G108), .ZN(G238) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U921 ( .A(n908), .B(n818), .ZN(n819) );
  NOR2_X1 U922 ( .A1(G860), .A2(n819), .ZN(n820) );
  XOR2_X1 U923 ( .A(KEYINPUT83), .B(n820), .Z(n821) );
  XOR2_X1 U924 ( .A(n822), .B(n821), .Z(G145) );
  XOR2_X1 U925 ( .A(G2100), .B(G2096), .Z(n824) );
  XNOR2_X1 U926 ( .A(KEYINPUT42), .B(G2678), .ZN(n823) );
  XNOR2_X1 U927 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2090), .Z(n826) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n825) );
  XNOR2_X1 U930 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U931 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2084), .ZN(n829) );
  XNOR2_X1 U933 ( .A(n830), .B(n829), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1976), .B(G1981), .Z(n832) );
  XNOR2_X1 U935 ( .A(G1986), .B(G1966), .ZN(n831) );
  XNOR2_X1 U936 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U937 ( .A(n833), .B(G2474), .Z(n835) );
  XNOR2_X1 U938 ( .A(G1956), .B(G1971), .ZN(n834) );
  XNOR2_X1 U939 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1961), .Z(n837) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U942 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G136), .A2(n866), .ZN(n841) );
  NAND2_X1 U945 ( .A1(G100), .A2(n867), .ZN(n840) );
  NAND2_X1 U946 ( .A1(n841), .A2(n840), .ZN(n846) );
  NAND2_X1 U947 ( .A1(G124), .A2(n872), .ZN(n842) );
  XNOR2_X1 U948 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U949 ( .A1(G112), .A2(n870), .ZN(n843) );
  NAND2_X1 U950 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U951 ( .A1(n846), .A2(n845), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G142), .A2(n866), .ZN(n848) );
  NAND2_X1 U953 ( .A1(G106), .A2(n867), .ZN(n847) );
  NAND2_X1 U954 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U955 ( .A(n849), .B(KEYINPUT45), .ZN(n851) );
  NAND2_X1 U956 ( .A1(G130), .A2(n872), .ZN(n850) );
  NAND2_X1 U957 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G118), .A2(n870), .ZN(n852) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(n852), .ZN(n853) );
  NOR2_X1 U960 ( .A1(n854), .A2(n853), .ZN(n858) );
  XOR2_X1 U961 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n856) );
  XNOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n855) );
  XNOR2_X1 U963 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U964 ( .A(n858), .B(n857), .ZN(n861) );
  XOR2_X1 U965 ( .A(G160), .B(n859), .Z(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n865) );
  XNOR2_X1 U967 ( .A(G162), .B(n862), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n863), .B(n936), .ZN(n864) );
  XOR2_X1 U969 ( .A(n865), .B(n864), .Z(n880) );
  NAND2_X1 U970 ( .A1(G139), .A2(n866), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G103), .A2(n867), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G115), .A2(n870), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(KEYINPUT112), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G127), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT113), .B(n878), .Z(n931) );
  XNOR2_X1 U980 ( .A(G164), .B(n931), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U982 ( .A(n882), .B(n881), .Z(n883) );
  NOR2_X1 U983 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U984 ( .A(G171), .B(G286), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(n886), .B(n917), .Z(n887) );
  NOR2_X1 U987 ( .A1(G37), .A2(n887), .ZN(G397) );
  XOR2_X1 U988 ( .A(G2443), .B(G2427), .Z(n889) );
  XNOR2_X1 U989 ( .A(G2438), .B(G2454), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(n890), .B(G2435), .Z(n892) );
  XNOR2_X1 U992 ( .A(G1341), .B(G1348), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U994 ( .A(G2430), .B(G2446), .Z(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT106), .B(G2451), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U997 ( .A(n896), .B(n895), .Z(n897) );
  NAND2_X1 U998 ( .A1(G14), .A2(n897), .ZN(n903) );
  NAND2_X1 U999 ( .A1(n903), .A2(G319), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n898), .ZN(n899) );
  NOR2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(n903), .ZN(G401) );
  XNOR2_X1 U1007 ( .A(KEYINPUT56), .B(G16), .ZN(n929) );
  XNOR2_X1 U1008 ( .A(G1966), .B(G168), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(n906), .B(KEYINPUT57), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n907), .B(G1956), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n908), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(G301), .B(G1961), .ZN(n909) );
  NOR2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(G1348), .B(n917), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n927) );
  XNOR2_X1 U1020 ( .A(G1971), .B(G303), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT121), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT122), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(KEYINPUT123), .ZN(n1011) );
  XNOR2_X1 U1028 ( .A(G2072), .B(n931), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G164), .B(G2078), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(n932), .B(KEYINPUT118), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT50), .ZN(n954) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G160), .ZN(n949) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT116), .B(n940), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n943), .Z(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT117), .B(n950), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1046 ( .A(KEYINPUT52), .B(n955), .Z(n956) );
  NOR2_X1 U1047 ( .A1(KEYINPUT55), .A2(n956), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT119), .B(n957), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n958), .A2(G29), .ZN(n1009) );
  XOR2_X1 U1050 ( .A(n959), .B(G27), .Z(n962) );
  XOR2_X1 U1051 ( .A(n960), .B(G32), .Z(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n970) );
  XOR2_X1 U1053 ( .A(G25), .B(G1991), .Z(n963) );
  NAND2_X1 U1054 ( .A1(n963), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G26), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G2072), .B(G33), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1058 ( .A(KEYINPUT120), .B(n966), .Z(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(KEYINPUT53), .ZN(n974) );
  XOR2_X1 U1062 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G35), .B(G2090), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT55), .B(n977), .Z(n978) );
  NOR2_X1 U1068 ( .A1(G29), .A2(n978), .ZN(n1007) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G23), .B(G1976), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1072 ( .A(G1986), .B(G24), .Z(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  XOR2_X1 U1074 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n983) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n999) );
  XOR2_X1 U1076 ( .A(G1966), .B(G21), .Z(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n985), .ZN(n997) );
  XNOR2_X1 U1078 ( .A(G20), .B(n986), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G1981), .B(G6), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT59), .B(G1348), .Z(n991) );
  XNOR2_X1 U1084 ( .A(G4), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT124), .B(n994), .Z(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT60), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G5), .B(G1961), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT61), .B(n1002), .ZN(n1004) );
  INV_X1 U1093 ( .A(G16), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(G11), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1012), .Z(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1013), .ZN(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

