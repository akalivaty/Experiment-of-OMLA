//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n469), .B2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n461), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n461), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n461), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n482), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n500), .A2(KEYINPUT68), .A3(new_n491), .A4(new_n490), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(G50), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G166));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n514), .A2(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT70), .B(G51), .Z(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT69), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n524), .A2(new_n526), .A3(new_n529), .A4(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(new_n521), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n531), .A2(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n523), .A2(new_n530), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n522), .A2(G90), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n520), .B2(new_n521), .ZN(new_n542));
  AND2_X1   g117(.A1(G77), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n526), .A2(new_n529), .A3(G52), .A4(G543), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n507), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n526), .A2(new_n529), .A3(G43), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(KEYINPUT73), .B2(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n526), .A2(new_n529), .A3(G543), .A4(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n507), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n522), .B2(G91), .ZN(new_n572));
  INV_X1    g147(.A(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n516), .B2(KEYINPUT69), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n567), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n574), .A2(new_n526), .A3(new_n575), .A4(new_n564), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n568), .A2(new_n572), .A3(new_n576), .ZN(G299));
  XOR2_X1   g152(.A(new_n518), .B(KEYINPUT74), .Z(G303));
  AND3_X1   g153(.A1(new_n526), .A2(new_n529), .A3(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n522), .A2(G87), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(G651), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n505), .B2(new_n506), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(G73), .B2(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n531), .A2(KEYINPUT75), .A3(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n531), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(G48), .A2(G543), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(new_n514), .B2(new_n515), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n579), .A2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n516), .A2(new_n531), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT76), .B(G85), .Z(new_n598));
  OAI221_X1 g173(.A(new_n595), .B1(new_n584), .B2(new_n596), .C1(new_n597), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(KEYINPUT77), .A2(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(KEYINPUT77), .A2(KEYINPUT10), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n602), .A2(KEYINPUT78), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  INV_X1    g180(.A(new_n603), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n601), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n597), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n522), .A2(G92), .A3(new_n607), .A4(new_n604), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n520), .B2(new_n521), .ZN(new_n614));
  AND2_X1   g189(.A1(G79), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n526), .A2(new_n529), .A3(G54), .A4(G543), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT79), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n612), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n600), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n600), .B1(new_n622), .B2(G868), .ZN(G321));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G299), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(G168), .ZN(G297));
  XNOR2_X1  g202(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n464), .A2(new_n462), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  AOI22_X1  g215(.A1(G123), .A2(new_n482), .B1(new_n480), .B2(G135), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n461), .A2(KEYINPUT81), .A3(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(KEYINPUT81), .B1(new_n461), .B2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n648), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(KEYINPUT83), .A3(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n656), .B(new_n659), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n667), .B2(new_n662), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n664), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n673), .B(KEYINPUT17), .Z(new_n680));
  INV_X1    g255(.A(new_n671), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n676), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n673), .A3(new_n671), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n681), .A3(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(new_n697), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n693), .A2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n700), .A2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n706), .B1(new_n703), .B2(new_n704), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n709), .B1(new_n707), .B2(new_n710), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n690), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n715), .A2(new_n689), .A3(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G33), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G139), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n465), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n461), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT98), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n720), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2072), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G160), .B2(new_n719), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n719), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n719), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT29), .Z(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G2084), .B2(new_n736), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n740), .B2(new_n741), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n731), .A2(new_n737), .A3(new_n743), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n744), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1956), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n622), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n719), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G128), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(new_n719), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  NOR2_X1   g344(.A1(G171), .A2(new_n744), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G5), .B2(new_n744), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n482), .A2(G129), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n462), .A2(G105), .ZN(new_n778));
  INV_X1    g353(.A(G141), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n465), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n719), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n719), .B2(G32), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT30), .B(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(new_n719), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n645), .B2(new_n719), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n772), .B(new_n791), .C1(new_n783), .C2(new_n784), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n555), .B2(G16), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(G1341), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G1341), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n771), .B2(new_n769), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n792), .A2(new_n795), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n750), .A2(new_n754), .A3(new_n758), .A4(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT99), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n744), .A2(G6), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n593), .B2(new_n744), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT92), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n581), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G49), .B2(new_n579), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n744), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n744), .B2(G23), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n744), .A2(G22), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G166), .B2(new_n744), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1971), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n808), .A2(new_n809), .A3(new_n816), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  MUX2_X1   g400(.A(G24), .B(G290), .S(G16), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1986), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n719), .A2(G25), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT89), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n482), .A2(G119), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT90), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G107), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n480), .B2(G131), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n829), .B1(new_n836), .B2(G29), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G1991), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n827), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n824), .A2(new_n825), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n824), .A2(new_n825), .A3(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT94), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(KEYINPUT36), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT96), .B(KEYINPUT36), .Z(new_n848));
  AOI22_X1  g423(.A1(new_n846), .A2(new_n847), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n843), .A2(KEYINPUT95), .A3(KEYINPUT36), .A4(new_n845), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n803), .B1(new_n849), .B2(new_n850), .ZN(G311));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n803), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(G150));
  NAND2_X1  g429(.A1(new_n622), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT38), .Z(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n507), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G651), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n526), .A2(new_n529), .A3(G55), .A4(G543), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n522), .A2(G93), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n554), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n554), .A2(new_n863), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n856), .B(new_n866), .Z(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  XNOR2_X1  g448(.A(new_n781), .B(new_n765), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n497), .A2(KEYINPUT100), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n500), .A2(new_n876), .A3(new_n491), .A4(new_n490), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(KEYINPUT101), .B2(new_n728), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n728), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n729), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n878), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n874), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n836), .B(new_n636), .Z(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  INV_X1    g463(.A(G118), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G130), .B2(new_n482), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n480), .A2(G142), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n836), .B(new_n636), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n896), .A2(KEYINPUT103), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT103), .B1(new_n896), .B2(new_n899), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n880), .B(new_n886), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n886), .A2(new_n880), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n896), .A2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n897), .B(new_n895), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT103), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n645), .B(G162), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G160), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n909), .B(new_n914), .C1(new_n903), .C2(new_n904), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g492(.A(new_n631), .B(new_n866), .ZN(new_n918));
  NAND2_X1  g493(.A1(G299), .A2(KEYINPUT104), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n568), .A2(new_n572), .A3(new_n576), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n622), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT79), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT79), .B1(new_n616), .B2(new_n617), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n611), .B(new_n610), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(KEYINPUT104), .A3(G299), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n918), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n811), .A2(KEYINPUT105), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NOR2_X1   g512(.A1(G288), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n593), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n811), .A2(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g515(.A1(G288), .A2(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G305), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(G166), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G290), .B(new_n518), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n939), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n935), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n935), .A2(new_n949), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n625), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n863), .A2(new_n625), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(G295));
  INV_X1    g530(.A(new_n954), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT106), .ZN(G331));
  AND2_X1   g533(.A1(G286), .A2(G301), .ZN(new_n959));
  NOR2_X1   g534(.A1(G286), .A2(G301), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n864), .A2(new_n865), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G168), .A2(G171), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n550), .A2(G651), .B1(new_n522), .B2(G81), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n859), .A2(G651), .B1(new_n522), .B2(G93), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n552), .A4(new_n861), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n554), .A2(new_n863), .ZN(new_n966));
  NAND2_X1  g541(.A1(G286), .A2(G301), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n962), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n968), .A3(KEYINPUT108), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n866), .A2(new_n970), .A3(new_n967), .A4(new_n962), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n961), .A2(new_n968), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n933), .A2(new_n972), .B1(new_n927), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n974), .B2(new_n949), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n927), .B1(new_n969), .B2(new_n971), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT41), .B1(new_n922), .B2(new_n926), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n981), .B2(new_n973), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(new_n948), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n931), .A2(new_n932), .A3(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n972), .A2(new_n928), .ZN(new_n985));
  AND4_X1   g560(.A1(new_n977), .A2(new_n948), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n975), .B(new_n976), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n985), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT109), .B1(new_n990), .B2(new_n949), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n982), .A2(new_n977), .A3(new_n948), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .A3(new_n976), .A4(new_n975), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n990), .B2(new_n949), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n983), .B2(new_n986), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n993), .A2(new_n975), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT44), .B1(new_n1002), .B2(new_n976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(new_n781), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n884), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n480), .A2(G137), .B1(G101), .B2(new_n462), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n475), .B1(new_n474), .B2(G2105), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT67), .B(new_n461), .C1(new_n472), .C2(new_n473), .ZN(new_n1013));
  OAI211_X1 g588(.A(G40), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1008), .A2(KEYINPUT111), .A3(new_n1009), .A4(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(G1996), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1005), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2067), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n765), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n1019), .B2(new_n781), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1018), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n836), .B(new_n838), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G290), .B(G1986), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1018), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n580), .A2(G1976), .A3(new_n581), .A4(new_n582), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n497), .A2(new_n1007), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1034), .B(G8), .C1(new_n1014), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n811), .A2(G1976), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1037), .A2(new_n1033), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n587), .A2(new_n588), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G651), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  INV_X1    g621(.A(new_n592), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n589), .B2(new_n592), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT49), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1014), .B2(new_n1035), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT117), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1053), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n1055), .A2(new_n1050), .A3(new_n1056), .A4(new_n1051), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1042), .B(new_n1043), .C1(new_n1054), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G303), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT55), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n502), .B2(new_n1007), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(G160), .B(G40), .C1(new_n1035), .C2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1064), .A2(new_n1067), .A3(G2090), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n502), .A2(new_n1007), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT113), .A3(new_n1009), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n1007), .A4(new_n877), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(new_n1016), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1384), .B1(new_n499), .B2(new_n501), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(KEYINPUT45), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1971), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(KEYINPUT114), .A3(new_n1077), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1060), .B(new_n1062), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1014), .B1(new_n1009), .B2(new_n1035), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1069), .B2(new_n1009), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n747), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n497), .A2(new_n1007), .A3(new_n1065), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n1014), .ZN(new_n1087));
  INV_X1    g662(.A(G2084), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1087), .B(new_n1088), .C1(new_n1063), .C2(new_n1074), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(G8), .A4(G168), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1074), .A2(new_n1063), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1014), .B1(new_n1035), .B2(new_n1066), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G2090), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1092), .B1(new_n1098), .B2(new_n1062), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1059), .B1(new_n1082), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1062), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1068), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1081), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1104), .B2(G8), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1088), .A2(new_n1106), .B1(new_n1084), .B2(new_n747), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1107), .A2(new_n1060), .A3(G286), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1059), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT63), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1111), .A2(G1976), .A3(G288), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n589), .A2(G1981), .A3(new_n592), .ZN(new_n1113));
  OAI221_X1 g688(.A(G8), .B1(new_n1014), .B2(new_n1035), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1100), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1087), .B(KEYINPUT118), .C1(new_n1063), .C2(new_n1074), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n757), .A3(new_n1119), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1014), .A2(G2067), .A3(new_n1035), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1070), .A2(new_n1072), .A3(new_n1075), .A4(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(G299), .B(KEYINPUT57), .Z(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1096), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n622), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1128), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1070), .A2(new_n1072), .A3(new_n1075), .A4(new_n1019), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1014), .B2(new_n1035), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1139), .B2(new_n555), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n554), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1124), .A2(new_n1127), .A3(new_n1125), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1125), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n925), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n925), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT60), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1133), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n1162));
  NAND2_X1  g737(.A1(G286), .A2(G8), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT121), .Z(new_n1164));
  OAI211_X1 g739(.A(new_n1162), .B(new_n1164), .C1(new_n1107), .C2(new_n1060), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT51), .B1(new_n1107), .B2(new_n1164), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1164), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1090), .B2(G8), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1076), .B2(G2078), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1118), .A2(new_n769), .A3(new_n1119), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1170), .A2(G2078), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1084), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(G171), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n468), .A2(new_n461), .ZN(new_n1177));
  INV_X1    g752(.A(G40), .ZN(new_n1178));
  NOR4_X1   g753(.A1(new_n1177), .A2(new_n467), .A3(new_n1178), .A4(new_n1173), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1010), .A2(new_n1071), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1171), .A2(G301), .A3(new_n1172), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1169), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1097), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1062), .B1(new_n1185), .B2(new_n1060), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1059), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1082), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1171), .A2(new_n1172), .A3(new_n1180), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1171), .A2(KEYINPUT122), .A3(new_n1172), .A4(new_n1180), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(G171), .A3(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1171), .A2(G301), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1194), .A2(KEYINPUT54), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1184), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1115), .B(new_n1116), .C1(new_n1161), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1169), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1176), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT62), .B(new_n1165), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1104), .A2(G8), .A3(new_n1101), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1205), .A2(new_n1186), .A3(new_n1059), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1199), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1203), .A2(new_n1202), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1208), .A2(new_n1188), .A3(KEYINPUT124), .A4(new_n1201), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1198), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1133), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1144), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n622), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n1154), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1158), .B1(new_n1220), .B2(new_n1153), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1212), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1184), .A2(new_n1196), .A3(new_n1188), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1116), .B1(new_n1224), .B2(new_n1115), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1032), .B1(new_n1211), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(new_n1026), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1018), .B1(new_n1005), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1020), .A2(KEYINPUT46), .A3(new_n1023), .ZN(new_n1229));
  AOI21_X1  g804(.A(KEYINPUT46), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT47), .ZN(new_n1232));
  OR2_X1    g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1235));
  AND3_X1   g810(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1234), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1237));
  AND3_X1   g812(.A1(new_n831), .A2(new_n838), .A3(new_n835), .ZN(new_n1238));
  AOI22_X1  g813(.A1(new_n1028), .A2(new_n1238), .B1(new_n1025), .B2(new_n766), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1022), .A2(G1986), .A3(G290), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1240), .B(KEYINPUT48), .ZN(new_n1241));
  OAI22_X1  g816(.A1(new_n1239), .A2(new_n1022), .B1(new_n1030), .B2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n1236), .A2(new_n1237), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1226), .A2(new_n1243), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g819(.A1(G227), .A2(new_n459), .ZN(new_n1246));
  NAND3_X1  g820(.A1(new_n669), .A2(new_n717), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g821(.A(new_n1247), .B1(new_n913), .B2(new_n915), .ZN(new_n1248));
  AND3_X1   g822(.A1(new_n998), .A2(new_n1248), .A3(KEYINPUT126), .ZN(new_n1249));
  AOI21_X1  g823(.A(KEYINPUT126), .B1(new_n998), .B2(new_n1248), .ZN(new_n1250));
  OAI21_X1  g824(.A(KEYINPUT127), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n998), .A2(new_n1248), .ZN(new_n1252));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1255));
  NAND3_X1  g829(.A1(new_n998), .A2(new_n1248), .A3(KEYINPUT126), .ZN(new_n1256));
  NAND3_X1  g830(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AND2_X1   g831(.A1(new_n1251), .A2(new_n1257), .ZN(G308));
  NAND2_X1  g832(.A1(new_n1254), .A2(new_n1256), .ZN(G225));
endmodule


