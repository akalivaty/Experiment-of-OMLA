//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n476), .A2(KEYINPUT4), .A3(G138), .ZN(new_n485));
  NAND2_X1  g060(.A1(G102), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n476), .B2(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n490), .B2(new_n462), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n476), .A2(G138), .A3(new_n462), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT5), .B(G543), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n495), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n494), .B(new_n496), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT71), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n497), .A2(new_n498), .A3(G651), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(new_n504), .B1(KEYINPUT6), .B2(new_n495), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(new_n494), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G88), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n494), .A2(G62), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n504), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n496), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n515), .B2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n508), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n505), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n494), .A2(G63), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G51), .B1(G651), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n521), .A3(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n494), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n523), .A2(G52), .B1(G651), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n502), .A2(new_n507), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n508), .A2(G81), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n494), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT72), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G43), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n537), .A2(new_n540), .A3(KEYINPUT73), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND4_X1  g127(.A1(new_n512), .A2(G53), .A3(G543), .A4(new_n496), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n505), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n502), .A2(G91), .A3(new_n507), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n494), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT74), .Z(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(G299));
  OR2_X1    g138(.A1(new_n494), .A2(G74), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n523), .A2(G49), .B1(G651), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n534), .ZN(G288));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n529), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n522), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n502), .A2(G86), .A3(new_n507), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n502), .A2(new_n507), .A3(KEYINPUT75), .A4(G86), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n529), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n523), .A2(G47), .B1(G651), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n534), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n523), .A2(G54), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OR2_X1    g165(.A1(KEYINPUT77), .A2(G66), .ZN(new_n591));
  NAND2_X1  g166(.A1(KEYINPUT77), .A2(G66), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n494), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n495), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n534), .B2(new_n598), .ZN(new_n599));
  AOI211_X1 g174(.A(new_n590), .B(new_n595), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n604), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(G868), .B2(new_n604), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n480), .A2(G2104), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT79), .B1(new_n480), .B2(G135), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G123), .B2(new_n478), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n480), .A2(KEYINPUT79), .A3(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n624), .ZN(G156));
  INV_X1    g200(.A(G14), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  OAI21_X1  g205(.A(KEYINPUT14), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n630), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(KEYINPUT82), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n641), .A2(new_n642), .A3(new_n647), .A4(new_n644), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n626), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n645), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT17), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n661), .C1(new_n659), .C2(new_n655), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(KEYINPUT20), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(KEYINPUT20), .C2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT83), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n678), .B(new_n683), .ZN(G229));
  NAND2_X1  g259(.A1(G171), .A2(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G5), .B2(G16), .ZN(new_n686));
  INV_X1    g261(.A(G1961), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n688));
  OR2_X1    g263(.A1(KEYINPUT24), .A2(G34), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(KEYINPUT24), .A2(G34), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G160), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G2084), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G2090), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(G29), .A2(G33), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n480), .A2(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n462), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n690), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n623), .A2(new_n690), .ZN(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n711), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n700), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n695), .B(new_n717), .C1(new_n688), .C2(new_n694), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n719));
  INV_X1    g294(.A(G26), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G29), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n723));
  INV_X1    g298(.A(G104), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n462), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT94), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n478), .A2(G128), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n480), .A2(G140), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n722), .B1(new_n729), .B2(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n719), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G2067), .ZN(new_n732));
  INV_X1    g307(.A(G32), .ZN(new_n733));
  AOI21_X1  g308(.A(KEYINPUT97), .B1(new_n690), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G141), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n478), .A2(G129), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n690), .ZN(new_n744));
  MUX2_X1   g319(.A(new_n734), .B(KEYINPUT97), .S(new_n744), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n693), .A2(G2084), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n731), .A2(G2067), .ZN(new_n749));
  AND4_X1   g324(.A1(new_n732), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G11), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n718), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n690), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n690), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G2078), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n600), .B2(new_n756), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(G16), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI22_X1  g338(.A1(G299), .A2(G16), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1956), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n756), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n756), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n686), .A2(new_n687), .B1(new_n754), .B2(G2078), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n766), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n752), .A2(new_n755), .A3(new_n759), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n761), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n546), .B2(new_n761), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT93), .B(G1341), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT34), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT91), .B(G1971), .ZN(new_n779));
  NAND2_X1  g354(.A1(G303), .A2(new_n761), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n762), .A2(G22), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n780), .A2(new_n781), .A3(new_n779), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n578), .A2(new_n756), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G6), .B2(new_n756), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n784), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G288), .A2(G16), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n756), .A2(G23), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n795));
  OAI21_X1  g370(.A(G1976), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n795), .ZN(new_n797));
  INV_X1    g372(.A(G1976), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n797), .A2(new_n798), .A3(new_n793), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n778), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n800), .A2(new_n787), .A3(new_n778), .A4(new_n788), .ZN(new_n802));
  AOI22_X1  g377(.A1(G119), .A2(new_n478), .B1(new_n480), .B2(G131), .ZN(new_n803));
  OR2_X1    g378(.A1(G95), .A2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT85), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n463), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n806), .B1(new_n805), .B2(new_n804), .C1(G107), .C2(new_n462), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT88), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT35), .B(G1991), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT87), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT86), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n810), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n761), .A2(G24), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n585), .B(KEYINPUT76), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n761), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT90), .B(G1986), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n802), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT92), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n802), .A2(new_n822), .A3(new_n814), .A4(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n801), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI211_X1 g401(.A(KEYINPUT36), .B(new_n801), .C1(new_n821), .C2(new_n823), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n773), .B(new_n777), .C1(new_n826), .C2(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  NAND2_X1  g404(.A1(new_n523), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n494), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n495), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n508), .B2(G93), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n600), .A2(G559), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n546), .A2(new_n834), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(new_n542), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n844), .B2(KEYINPUT101), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(KEYINPUT101), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n846), .B2(new_n847), .ZN(G145));
  XOR2_X1   g423(.A(new_n623), .B(G162), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n743), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n462), .B1(new_n852), .B2(new_n488), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT4), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n492), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n485), .A2(new_n486), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n462), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n729), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n478), .A2(G130), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n480), .A2(G142), .ZN(new_n861));
  NOR2_X1   g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n614), .B(new_n707), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n851), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n743), .A3(new_n868), .ZN(new_n873));
  XOR2_X1   g448(.A(G160), .B(new_n808), .Z(new_n874));
  AND3_X1   g449(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n850), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  INV_X1    g453(.A(new_n874), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n743), .B1(new_n872), .B2(new_n868), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n869), .A2(new_n851), .A3(new_n870), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n849), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g461(.A(new_n595), .B1(new_n596), .B2(new_n599), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n589), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n604), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(G299), .A3(new_n589), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n842), .A2(new_n607), .A3(new_n600), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n840), .A2(new_n609), .A3(new_n841), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(KEYINPUT102), .A3(new_n890), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n600), .A2(KEYINPUT102), .A3(G299), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n896), .A2(new_n897), .A3(new_n902), .A4(new_n898), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n893), .A2(new_n894), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  AOI211_X1 g483(.A(new_n908), .B(new_n895), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n816), .B(G288), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G290), .B(G288), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n578), .B(G303), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OR3_X1    g492(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n907), .A2(new_n909), .A3(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n833), .A2(G868), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G295));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(G331));
  XNOR2_X1  g503(.A(G286), .B(G301), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n840), .A2(new_n841), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G171), .B(G286), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n833), .B1(new_n544), .B2(new_n545), .ZN(new_n932));
  INV_X1    g507(.A(new_n841), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n904), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n934), .A2(KEYINPUT106), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n891), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n878), .B1(new_n941), .B2(new_n919), .ZN(new_n942));
  INV_X1    g517(.A(new_n919), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n896), .A2(new_n897), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT41), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n891), .A2(new_n898), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n939), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n930), .A2(new_n934), .A3(new_n891), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT108), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n943), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n942), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n904), .A2(new_n935), .B1(new_n939), .B2(new_n891), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n943), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n941), .A2(new_n919), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT43), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n942), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(G397));
  XOR2_X1   g542(.A(new_n729), .B(G2067), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT110), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n743), .B(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n808), .B(new_n812), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT111), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n855), .B2(new_n857), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n981), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n729), .A2(G2067), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n808), .A2(new_n812), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n982), .A2(new_n985), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n981), .B1(new_n969), .B2(new_n851), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n970), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT46), .Z(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n994));
  XNOR2_X1  g569(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT115), .B(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT116), .Z(new_n999));
  INV_X1    g574(.A(new_n979), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n976), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(G8), .C1(new_n798), .C2(G288), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1002), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n1002), .B2(KEYINPUT52), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n999), .A2(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(new_n492), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n852), .A2(new_n488), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G2105), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1010), .B2(KEYINPUT4), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1006), .B(new_n1007), .C1(new_n1011), .C2(new_n487), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n976), .A2(new_n1014), .A3(new_n1006), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT113), .B1(new_n976), .B2(new_n1006), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1016), .A2(new_n1020), .A3(new_n1021), .A4(new_n1000), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n979), .B1(KEYINPUT45), .B2(new_n976), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n978), .ZN(new_n1024));
  INV_X1    g599(.A(G1971), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n1000), .A3(new_n1012), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G2090), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1971), .B1(new_n1023), .B2(new_n978), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1028), .B(KEYINPUT55), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n573), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n574), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n576), .A2(new_n577), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  AND4_X1   g619(.A1(KEYINPUT117), .A2(new_n1043), .A3(new_n1044), .A4(new_n1040), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT117), .B1(new_n578), .B2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1001), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT49), .B(new_n1042), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1049), .A2(new_n1056), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1005), .B(new_n1039), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1016), .A2(new_n1020), .A3(new_n1000), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  INV_X1    g635(.A(G2078), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1023), .A2(new_n978), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1059), .A2(new_n687), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n979), .B1(new_n976), .B2(new_n977), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(KEYINPUT45), .B2(new_n976), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1065), .A2(new_n1060), .A3(G2078), .ZN(new_n1066));
  AOI21_X1  g641(.A(G301), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n769), .ZN(new_n1068));
  INV_X1    g643(.A(G2084), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1016), .A2(new_n1020), .A3(new_n1069), .A4(new_n1000), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(G168), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g648(.A(G168), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  OAI211_X1 g650(.A(G8), .B(new_n1071), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT62), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1058), .A2(new_n1067), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1001), .A2(G2067), .ZN(new_n1082));
  INV_X1    g657(.A(G1348), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1082), .B(new_n600), .C1(new_n1059), .C2(new_n1083), .ZN(new_n1084));
  NOR4_X1   g659(.A1(G164), .A2(KEYINPUT112), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1014), .B1(new_n976), .B2(new_n1006), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1000), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1082), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n888), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT60), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT126), .B1(new_n1093), .B2(KEYINPUT125), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(G1341), .Z(new_n1096));
  OAI22_X1  g671(.A1(new_n1024), .A2(G1996), .B1(new_n1050), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1094), .B1(new_n1097), .B2(new_n546), .ZN(new_n1098));
  AOI211_X1 g673(.A(KEYINPUT60), .B(new_n1082), .C1(new_n1059), .C2(new_n1083), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n600), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT121), .B(G1956), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1033), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G299), .B(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT56), .B(G2072), .Z(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT123), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1023), .A2(new_n978), .A3(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1102), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT61), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1104), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1102), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1093), .A2(KEYINPUT126), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1097), .A2(new_n546), .A3(new_n1094), .A4(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1092), .A2(new_n1100), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1109), .B1(new_n1091), .B2(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G301), .B(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1059), .A2(new_n687), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1062), .A2(new_n1060), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n978), .A2(G40), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n469), .A2(new_n473), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(KEYINPUT53), .A3(new_n1061), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1126), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1125), .B(new_n1133), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1058), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1005), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1051), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1030), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1052), .B(KEYINPUT119), .Z(new_n1139));
  OR2_X1    g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1081), .A2(new_n1135), .A3(new_n1138), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1072), .A2(G286), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1058), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1058), .A2(KEYINPUT120), .A3(new_n1145), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1137), .A2(new_n1030), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(new_n1149), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1136), .A2(new_n1031), .A3(new_n1145), .A4(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1144), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G290), .A2(G1986), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n975), .A2(new_n1156), .A3(new_n983), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(new_n980), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n996), .B1(new_n1155), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G227), .A2(new_n460), .ZN(new_n1161));
  INV_X1    g735(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(G229), .B1(new_n649), .B2(new_n650), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n885), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g738(.A(new_n955), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n1165), .A2(new_n956), .A3(new_n959), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n959), .A2(new_n960), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(KEYINPUT43), .ZN(new_n1168));
  AOI211_X1 g742(.A(new_n1162), .B(new_n1164), .C1(new_n1166), .C2(new_n1168), .ZN(G308));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n1170), .A2(new_n885), .A3(new_n1161), .A4(new_n1163), .ZN(G225));
endmodule


