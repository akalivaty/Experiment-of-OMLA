

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NAND2_X2 U556 ( .A1(n685), .A2(n787), .ZN(n731) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n526), .Z(n882) );
  NOR2_X1 U558 ( .A1(n689), .A2(n688), .ZN(n692) );
  OR2_X1 U559 ( .A1(n764), .A2(n763), .ZN(n520) );
  NOR2_X1 U560 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U561 ( .A(KEYINPUT29), .B(KEYINPUT103), .ZN(n712) );
  INV_X1 U562 ( .A(n978), .ZN(n748) );
  NOR2_X1 U563 ( .A1(n764), .A2(n748), .ZN(n749) );
  AND2_X1 U564 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U565 ( .A1(n765), .A2(n520), .ZN(n766) );
  OR2_X1 U566 ( .A1(n767), .A2(n766), .ZN(n806) );
  NOR2_X1 U567 ( .A1(G543), .A2(n542), .ZN(n539) );
  NOR2_X1 U568 ( .A1(G651), .A2(n649), .ZN(n655) );
  NOR2_X2 U569 ( .A1(G2105), .A2(n522), .ZN(n881) );
  XOR2_X1 U570 ( .A(KEYINPUT74), .B(n583), .Z(n972) );
  INV_X1 U571 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G101), .A2(n881), .ZN(n521) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n521), .Z(n525) );
  AND2_X1 U574 ( .A1(n522), .A2(G2105), .ZN(n877) );
  NAND2_X1 U575 ( .A1(G125), .A2(n877), .ZN(n523) );
  XOR2_X1 U576 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n882), .A2(G137), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U581 ( .A(KEYINPUT66), .B(n527), .Z(n878) );
  NAND2_X1 U582 ( .A1(G113), .A2(n878), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U584 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U585 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U586 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U587 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  INV_X1 U588 ( .A(G132), .ZN(G219) );
  NAND2_X1 U589 ( .A1(G69), .A2(G120), .ZN(n532) );
  NOR2_X1 U590 ( .A1(G237), .A2(n532), .ZN(n533) );
  NAND2_X1 U591 ( .A1(G108), .A2(n533), .ZN(n830) );
  NAND2_X1 U592 ( .A1(n830), .A2(G567), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G220), .A2(G219), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT22), .B(n534), .Z(n535) );
  NOR2_X1 U595 ( .A1(G218), .A2(n535), .ZN(n536) );
  NAND2_X1 U596 ( .A1(G96), .A2(n536), .ZN(n831) );
  NAND2_X1 U597 ( .A1(n831), .A2(G2106), .ZN(n537) );
  AND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(G319) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n658) );
  NAND2_X1 U600 ( .A1(G85), .A2(n658), .ZN(n541) );
  INV_X1 U601 ( .A(G651), .ZN(n542) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n539), .Z(n654) );
  NAND2_X1 U603 ( .A1(G60), .A2(n654), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n546) );
  XOR2_X1 U605 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  NOR2_X1 U606 ( .A1(n649), .A2(n542), .ZN(n652) );
  NAND2_X1 U607 ( .A1(G72), .A2(n652), .ZN(n544) );
  NAND2_X1 U608 ( .A1(G47), .A2(n655), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U610 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U611 ( .A1(G64), .A2(n654), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G52), .A2(n655), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n658), .A2(G90), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT67), .B(n549), .Z(n551) );
  NAND2_X1 U616 ( .A1(n652), .A2(G77), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G102), .A2(n881), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G138), .A2(n882), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G126), .A2(n877), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G114), .A2(n878), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(G164) );
  XOR2_X1 U628 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n562) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n826) );
  NAND2_X1 U632 ( .A1(n826), .A2(G567), .ZN(n563) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U634 ( .A1(G56), .A2(n654), .ZN(n564) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n564), .Z(n571) );
  NAND2_X1 U636 ( .A1(G81), .A2(n658), .ZN(n565) );
  XNOR2_X1 U637 ( .A(n565), .B(KEYINPUT12), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n566), .B(KEYINPUT72), .ZN(n568) );
  NAND2_X1 U639 ( .A1(G68), .A2(n652), .ZN(n567) );
  NAND2_X1 U640 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(n569), .Z(n570) );
  NOR2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n655), .A2(G43), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n973) );
  INV_X1 U645 ( .A(n973), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n574), .A2(G860), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  INV_X1 U648 ( .A(G868), .ZN(n606) );
  NOR2_X1 U649 ( .A1(G301), .A2(n606), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G54), .A2(n655), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G79), .A2(n652), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n654), .A2(G66), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U654 ( .A1(G92), .A2(n658), .ZN(n577) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n577), .ZN(n578) );
  NOR2_X1 U656 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n582), .B(KEYINPUT15), .ZN(n583) );
  NOR2_X1 U659 ( .A1(n972), .A2(G868), .ZN(n584) );
  NOR2_X1 U660 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n658), .A2(G89), .ZN(n586) );
  XNOR2_X1 U662 ( .A(n586), .B(KEYINPUT4), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G76), .A2(n652), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U665 ( .A(KEYINPUT5), .B(n589), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n654), .A2(G63), .ZN(n590) );
  XOR2_X1 U667 ( .A(KEYINPUT75), .B(n590), .Z(n592) );
  NAND2_X1 U668 ( .A1(n655), .A2(G51), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U670 ( .A(KEYINPUT6), .B(n593), .Z(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT7), .B(n596), .ZN(G168) );
  XOR2_X1 U673 ( .A(G168), .B(KEYINPUT8), .Z(n597) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n597), .ZN(G286) );
  NAND2_X1 U675 ( .A1(n652), .A2(G78), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT68), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G91), .A2(n658), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT69), .B(n601), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G65), .A2(n654), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G53), .A2(n655), .ZN(n602) );
  AND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(G299) );
  NAND2_X1 U684 ( .A1(G868), .A2(G286), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G299), .A2(n606), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U687 ( .A(G559), .ZN(n609) );
  NOR2_X1 U688 ( .A1(G860), .A2(n609), .ZN(n610) );
  XNOR2_X1 U689 ( .A(KEYINPUT77), .B(n610), .ZN(n611) );
  INV_X1 U690 ( .A(n972), .ZN(n633) );
  NAND2_X1 U691 ( .A1(n611), .A2(n633), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n973), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n633), .A2(G868), .ZN(n613) );
  NOR2_X1 U695 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G135), .A2(n882), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT78), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G123), .A2(n877), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G99), .A2(n881), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G111), .A2(n878), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n922) );
  XNOR2_X1 U706 ( .A(n922), .B(G2096), .ZN(n625) );
  INV_X1 U707 ( .A(G2100), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(G156) );
  NAND2_X1 U709 ( .A1(G80), .A2(n652), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G93), .A2(n658), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n654), .A2(G67), .ZN(n628) );
  XNOR2_X1 U713 ( .A(n628), .B(KEYINPUT80), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G55), .A2(n655), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n665) );
  NAND2_X1 U717 ( .A1(G559), .A2(n633), .ZN(n673) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n973), .Z(n634) );
  XNOR2_X1 U719 ( .A(n673), .B(n634), .ZN(n635) );
  NOR2_X1 U720 ( .A1(G860), .A2(n635), .ZN(n636) );
  XNOR2_X1 U721 ( .A(n665), .B(n636), .ZN(G145) );
  NAND2_X1 U722 ( .A1(G88), .A2(n658), .ZN(n637) );
  XNOR2_X1 U723 ( .A(n637), .B(KEYINPUT84), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G75), .A2(n652), .ZN(n639) );
  NAND2_X1 U725 ( .A1(G50), .A2(n655), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U727 ( .A1(G62), .A2(n654), .ZN(n640) );
  XNOR2_X1 U728 ( .A(KEYINPUT83), .B(n640), .ZN(n641) );
  NOR2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(G303) );
  INV_X1 U731 ( .A(G303), .ZN(G166) );
  NAND2_X1 U732 ( .A1(G49), .A2(n655), .ZN(n646) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n654), .A2(n647), .ZN(n648) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n648), .Z(n651) );
  NAND2_X1 U737 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G73), .A2(n652), .ZN(n653) );
  XNOR2_X1 U740 ( .A(n653), .B(KEYINPUT2), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G61), .A2(n654), .ZN(n657) );
  NAND2_X1 U742 ( .A1(G48), .A2(n655), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n658), .A2(G86), .ZN(n659) );
  XOR2_X1 U745 ( .A(KEYINPUT82), .B(n659), .Z(n660) );
  NOR2_X1 U746 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n663), .A2(n662), .ZN(G305) );
  NOR2_X1 U748 ( .A1(n665), .A2(G868), .ZN(n664) );
  XNOR2_X1 U749 ( .A(KEYINPUT87), .B(n664), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n665), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n666), .B(KEYINPUT85), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n667), .B(G290), .ZN(n670) );
  XNOR2_X1 U753 ( .A(G299), .B(n973), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U755 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U756 ( .A(G166), .B(n671), .ZN(n672) );
  XNOR2_X1 U757 ( .A(n672), .B(G305), .ZN(n894) );
  XNOR2_X1 U758 ( .A(n894), .B(n673), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(G868), .ZN(n675) );
  XNOR2_X1 U760 ( .A(KEYINPUT86), .B(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n681), .A2(G2072), .ZN(G158) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT88), .B(n682), .Z(n683) );
  NAND2_X1 U769 ( .A1(n683), .A2(G319), .ZN(n684) );
  XNOR2_X1 U770 ( .A(n684), .B(KEYINPUT89), .ZN(n829) );
  NAND2_X1 U771 ( .A1(n829), .A2(G36), .ZN(G176) );
  XOR2_X1 U772 ( .A(KEYINPUT27), .B(KEYINPUT101), .Z(n687) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n788) );
  INV_X1 U774 ( .A(n788), .ZN(n685) );
  XNOR2_X2 U775 ( .A(KEYINPUT99), .B(n731), .ZN(n715) );
  NAND2_X1 U776 ( .A1(G2072), .A2(n715), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n687), .B(n686), .ZN(n689) );
  INV_X1 U778 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U779 ( .A1(n715), .A2(n1006), .ZN(n688) );
  INV_X1 U780 ( .A(G299), .ZN(n983) );
  NOR2_X1 U781 ( .A1(n692), .A2(n983), .ZN(n691) );
  XOR2_X1 U782 ( .A(KEYINPUT28), .B(KEYINPUT102), .Z(n690) );
  XNOR2_X1 U783 ( .A(n691), .B(n690), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n983), .A2(n692), .ZN(n709) );
  XNOR2_X1 U785 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n699) );
  NOR2_X1 U786 ( .A1(G1996), .A2(n699), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n693), .A2(n973), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n715), .ZN(n695) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n731), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n972), .A2(n705), .ZN(n696) );
  NAND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n704) );
  INV_X1 U793 ( .A(G1341), .ZN(n1007) );
  NAND2_X1 U794 ( .A1(n1007), .A2(n699), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n698), .A2(n731), .ZN(n702) );
  INV_X1 U796 ( .A(G1996), .ZN(n808) );
  NOR2_X1 U797 ( .A1(n731), .A2(n808), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n972), .A2(n705), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n713), .B(n712), .ZN(n720) );
  INV_X1 U805 ( .A(G1961), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n714), .A2(n731), .ZN(n717) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .ZN(n950) );
  NAND2_X1 U808 ( .A1(n715), .A2(n950), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n725) );
  AND2_X1 U810 ( .A1(n725), .A2(G171), .ZN(n718) );
  XOR2_X1 U811 ( .A(KEYINPUT100), .B(n718), .Z(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n730) );
  NAND2_X1 U813 ( .A1(G8), .A2(n731), .ZN(n764) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n764), .ZN(n742) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n731), .ZN(n739) );
  NOR2_X1 U816 ( .A1(n742), .A2(n739), .ZN(n721) );
  NAND2_X1 U817 ( .A1(G8), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U820 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U821 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n728), .Z(n729) );
  NAND2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n740), .A2(G286), .ZN(n736) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n764), .ZN(n733) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n734), .A2(G303), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n737), .A2(G8), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n738), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U833 ( .A1(G8), .A2(n739), .ZN(n744) );
  INV_X1 U834 ( .A(n740), .ZN(n741) );
  NOR2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n760) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n754), .A2(n747), .ZN(n979) );
  NAND2_X1 U841 ( .A1(n760), .A2(n979), .ZN(n750) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n751), .ZN(n752) );
  XNOR2_X1 U844 ( .A(n752), .B(KEYINPUT105), .ZN(n753) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n969) );
  NAND2_X1 U846 ( .A1(n753), .A2(n969), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U848 ( .A1(n755), .A2(n764), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U851 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n764), .A2(n761), .ZN(n765) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U855 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NAND2_X1 U856 ( .A1(G119), .A2(n877), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G107), .A2(n878), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT95), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G95), .A2(n881), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n882), .A2(G131), .ZN(n773) );
  XOR2_X1 U863 ( .A(KEYINPUT96), .B(n773), .Z(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT97), .B(n776), .Z(n872) );
  INV_X1 U866 ( .A(G1991), .ZN(n948) );
  NOR2_X1 U867 ( .A1(n872), .A2(n948), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G129), .A2(n877), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G141), .A2(n882), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n878), .A2(G117), .ZN(n779) );
  XNOR2_X1 U872 ( .A(n779), .B(KEYINPUT98), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G105), .A2(n881), .ZN(n780) );
  XNOR2_X1 U874 ( .A(n780), .B(KEYINPUT38), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n888) );
  NOR2_X1 U877 ( .A1(n888), .A2(n808), .ZN(n785) );
  NOR2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n811) );
  XOR2_X1 U879 ( .A(G1986), .B(G290), .Z(n987) );
  NAND2_X1 U880 ( .A1(n811), .A2(n987), .ZN(n789) );
  NOR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n822) );
  NAND2_X1 U882 ( .A1(n789), .A2(n822), .ZN(n804) );
  XOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .Z(n821) );
  XNOR2_X1 U884 ( .A(KEYINPUT36), .B(KEYINPUT92), .ZN(n802) );
  NAND2_X1 U885 ( .A1(n882), .A2(G140), .ZN(n790) );
  XNOR2_X1 U886 ( .A(n790), .B(KEYINPUT90), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G104), .A2(n881), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n793), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n877), .A2(G128), .ZN(n794) );
  XOR2_X1 U891 ( .A(KEYINPUT91), .B(n794), .Z(n796) );
  NAND2_X1 U892 ( .A1(G116), .A2(n878), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U894 ( .A(n797), .B(KEYINPUT35), .Z(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U896 ( .A(KEYINPUT93), .B(n800), .Z(n801) );
  XOR2_X1 U897 ( .A(n802), .B(n801), .Z(n871) );
  AND2_X1 U898 ( .A1(n821), .A2(n871), .ZN(n803) );
  XNOR2_X1 U899 ( .A(n803), .B(KEYINPUT94), .ZN(n921) );
  NAND2_X1 U900 ( .A1(n921), .A2(n822), .ZN(n807) );
  AND2_X1 U901 ( .A1(n804), .A2(n807), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n820) );
  INV_X1 U903 ( .A(n807), .ZN(n818) );
  AND2_X1 U904 ( .A1(n808), .A2(n888), .ZN(n931) );
  AND2_X1 U905 ( .A1(n948), .A2(n872), .ZN(n923) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  XNOR2_X1 U907 ( .A(KEYINPUT106), .B(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n923), .A2(n810), .ZN(n812) );
  INV_X1 U909 ( .A(n811), .ZN(n928) );
  NOR2_X1 U910 ( .A1(n812), .A2(n928), .ZN(n813) );
  XOR2_X1 U911 ( .A(KEYINPUT107), .B(n813), .Z(n814) );
  NOR2_X1 U912 ( .A1(n931), .A2(n814), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT39), .B(n815), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n816), .A2(n822), .ZN(n817) );
  OR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  AND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n824) );
  NOR2_X1 U917 ( .A1(n821), .A2(n871), .ZN(n936) );
  NAND2_X1 U918 ( .A1(n936), .A2(n822), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(G2678), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U935 ( .A(KEYINPUT112), .B(G2090), .Z(n835) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2096), .B(G2100), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U941 ( .A(G2078), .B(G2084), .Z(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1986), .B(G1976), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1981), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G1991), .B(G1961), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1996), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT113), .B(G2474), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U952 ( .A(KEYINPUT41), .B(n850), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n851), .B(n1006), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G100), .A2(n881), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G136), .A2(n882), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n878), .A2(G112), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n854), .B(KEYINPUT114), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G124), .A2(n877), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n855), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n869) );
  NAND2_X1 U964 ( .A1(G127), .A2(n877), .ZN(n861) );
  NAND2_X1 U965 ( .A1(G115), .A2(n878), .ZN(n860) );
  NAND2_X1 U966 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n862), .B(KEYINPUT47), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G139), .A2(n882), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n881), .A2(G103), .ZN(n865) );
  XOR2_X1 U971 ( .A(KEYINPUT116), .B(n865), .Z(n866) );
  NOR2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n916) );
  XNOR2_X1 U973 ( .A(n916), .B(KEYINPUT48), .ZN(n868) );
  XNOR2_X1 U974 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U975 ( .A(G164), .B(n870), .ZN(n876) );
  XOR2_X1 U976 ( .A(n922), .B(G162), .Z(n874) );
  XOR2_X1 U977 ( .A(n872), .B(n871), .Z(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n892) );
  NAND2_X1 U980 ( .A1(G130), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n889) );
  XOR2_X1 U988 ( .A(n889), .B(n888), .Z(n890) );
  XNOR2_X1 U989 ( .A(G160), .B(n890), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G171), .B(G286), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n896), .B(n972), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2451), .B(G2443), .Z(n899) );
  XNOR2_X1 U997 ( .A(KEYINPUT109), .B(G2446), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT110), .B(G2438), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G2435), .B(G2454), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1002 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G2427), .B(KEYINPUT108), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G2430), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(n1007), .ZN(n907) );
  XOR2_X1 U1007 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1008 ( .A1(G14), .A2(n909), .ZN(n915) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n915), .ZN(G401) );
  INV_X1 U1018 ( .A(KEYINPUT55), .ZN(n964) );
  XOR2_X1 U1019 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1022 ( .A(KEYINPUT50), .B(n919), .Z(n939) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1026 ( .A(KEYINPUT117), .B(n924), .Z(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n929), .ZN(n934) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT119), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT52), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(n941), .B(KEYINPUT120), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n964), .A2(n942), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n943), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1041 ( .A(G2084), .B(G34), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT54), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n962) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n960) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n947), .B(G33), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(G25), .B(n948), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n949), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G27), .B(n950), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n960), .B(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n964), .B(n963), .ZN(n966) );
  INV_X1 U1060 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n967), .ZN(n1024) );
  INV_X1 U1063 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1064 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(n1020), .B(n968), .ZN(n994) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT57), .ZN(n992) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n972), .B(G1348), .ZN(n975) );
  XOR2_X1 U1071 ( .A(n1007), .B(n973), .Z(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n990) );
  AND2_X1 U1074 ( .A1(G303), .A2(G1971), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT124), .B(n982), .Z(n985) );
  XOR2_X1 U1078 ( .A(n983), .B(G1956), .Z(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT125), .B(n988), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1022) );
  XOR2_X1 U1085 ( .A(G1986), .B(G24), .Z(n998) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G23), .B(G1976), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n1000), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G5), .B(G1961), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .Z(n1005) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1005), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(n1006), .B(G20), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1007), .B(G19), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(G6), .B(G1981), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1012), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1015), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

