//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(KEYINPUT3), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G2104), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n462), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n462), .A2(new_n467), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n483), .A2(new_n468), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n486), .A2(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n468), .A3(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n477), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n468), .A2(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n462), .A2(new_n467), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n462), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT72), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT71), .B(G651), .Z(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT71), .B(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(new_n508), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n513), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n524), .A3(new_n513), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n512), .B1(new_n526), .B2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n523), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n523), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(G90), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n509), .A2(G64), .ZN(new_n540));
  AND2_X1   g115(.A1(G77), .A2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n515), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT74), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n523), .A2(G43), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n509), .A2(G56), .ZN(new_n549));
  AND2_X1   g124(.A1(G68), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n515), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n514), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT6), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n511), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n554), .A2(G81), .A3(new_n509), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n548), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT76), .B(G65), .Z(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n519), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n520), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n554), .A2(G53), .A3(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n523), .A2(new_n569), .A3(G53), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n568), .B1(new_n567), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n565), .B1(new_n572), .B2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  AND3_X1   g150(.A1(new_n521), .A2(new_n524), .A3(new_n513), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n576), .A2(new_n525), .B1(new_n510), .B2(new_n511), .ZN(G303));
  NAND2_X1  g152(.A1(G49), .A2(G543), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n516), .A2(KEYINPUT77), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n516), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n509), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n520), .A2(G87), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND4_X1  g159(.A1(new_n554), .A2(KEYINPUT80), .A3(G86), .A4(new_n509), .ZN(new_n585));
  OR2_X1    g160(.A1(KEYINPUT71), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(KEYINPUT71), .A2(G651), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n553), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n509), .B(G86), .C1(new_n588), .C2(new_n514), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n554), .A2(G48), .A3(G543), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n585), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  OAI21_X1  g170(.A(G61), .B1(new_n517), .B2(new_n518), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI211_X1 g172(.A(new_n595), .B(new_n511), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT78), .B1(new_n599), .B2(new_n515), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n507), .B2(new_n508), .ZN(new_n603));
  INV_X1    g178(.A(new_n597), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n515), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n599), .A2(KEYINPUT78), .A3(new_n515), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT79), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n593), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(G305));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n507), .B2(new_n508), .ZN(new_n614));
  AND2_X1   g189(.A1(G72), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n515), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n554), .A2(G85), .A3(new_n509), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n554), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G47), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n617), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n619), .B(KEYINPUT83), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n618), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n616), .B(KEYINPUT82), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G290));
  NAND2_X1  g206(.A1(new_n520), .A2(G92), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(G79), .A2(G543), .ZN(new_n637));
  INV_X1    g212(.A(G66), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n519), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n523), .A2(G54), .B1(new_n639), .B2(G651), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G868), .B2(G171), .ZN(G284));
  XOR2_X1   g218(.A(G284), .B(KEYINPUT85), .Z(G321));
  NAND2_X1  g219(.A1(G286), .A2(G868), .ZN(new_n645));
  INV_X1    g220(.A(new_n565), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n569), .B1(new_n523), .B2(G53), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT75), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n649), .B2(new_n571), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n650), .B2(G868), .ZN(G297));
  OAI21_X1  g226(.A(new_n645), .B1(new_n650), .B2(G868), .ZN(G280));
  INV_X1    g227(.A(new_n641), .ZN(new_n653));
  INV_X1    g228(.A(G559), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(G860), .ZN(G148));
  INV_X1    g230(.A(new_n556), .ZN(new_n656));
  INV_X1    g231(.A(G868), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n641), .A2(G559), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(new_n657), .ZN(G323));
  XNOR2_X1  g235(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g236(.A1(new_n484), .A2(G135), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  OR2_X1    g238(.A1(G99), .A2(G2105), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n664), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n665));
  INV_X1    g240(.A(G123), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n490), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(G2096), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT3), .B(G2104), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n470), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT13), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n670), .A2(new_n671), .A3(new_n678), .ZN(G156));
  XNOR2_X1  g254(.A(G2427), .B(G2438), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2430), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT15), .B(G2435), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(KEYINPUT14), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1341), .B(G1348), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2443), .B(G2446), .Z(new_n691));
  XNOR2_X1  g266(.A(G2451), .B(G2454), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(G14), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n694), .B2(new_n690), .ZN(G401));
  XOR2_X1   g271(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G2084), .B(G2090), .Z(new_n699));
  XNOR2_X1  g274(.A(G2067), .B(G2678), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT17), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G2072), .B(G2078), .Z(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n701), .B2(new_n697), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G2096), .B(G2100), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G227));
  XNOR2_X1  g284(.A(G1971), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT19), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1956), .B(G2474), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  XOR2_X1   g289(.A(G1961), .B(G1966), .Z(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT20), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n714), .A2(new_n715), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n720), .C1(new_n711), .C2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n721), .B(KEYINPUT92), .ZN(new_n726));
  INV_X1    g301(.A(new_n724), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(G1991), .B(G1996), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(G1981), .B(G1986), .ZN(new_n732));
  INV_X1    g307(.A(new_n730), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n725), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n731), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(G229));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n738), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2090), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n484), .A2(G139), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT25), .Z(new_n749));
  AOI22_X1  g324(.A1(new_n672), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n749), .C1(new_n468), .C2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n484), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n489), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(G105), .A2(new_n470), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n762), .A2(KEYINPUT96), .A3(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n738), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G32), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n738), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2084), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n753), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n744), .B(new_n746), .C1(new_n777), .C2(KEYINPUT97), .ZN(new_n778));
  INV_X1    g353(.A(G16), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G4), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n641), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n779), .A2(G21), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G286), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1966), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G11), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT31), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT31), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G28), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n738), .B1(new_n791), .B2(G28), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n668), .B2(G29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n785), .A2(new_n786), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n783), .A2(new_n787), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n753), .A2(KEYINPUT97), .A3(new_n770), .A4(new_n776), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n779), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n779), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT94), .B(G16), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(G19), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n556), .B2(new_n804), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1341), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n738), .A2(G26), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT28), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n484), .A2(G140), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n489), .A2(G128), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n468), .A2(G116), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G2067), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n738), .A2(G27), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G164), .B2(new_n738), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2078), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n807), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n798), .A2(new_n799), .A3(new_n802), .A4(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n801), .A2(G1961), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n767), .A2(new_n769), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n775), .A2(G2084), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n803), .A2(G20), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT23), .Z(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G299), .B2(G16), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1956), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n824), .A2(KEYINPUT98), .A3(new_n825), .A4(new_n826), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n778), .A2(new_n823), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n626), .A2(new_n630), .A3(new_n804), .ZN(new_n837));
  INV_X1    g412(.A(G1986), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n804), .A2(G24), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n484), .A2(G131), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n489), .A2(G119), .ZN(new_n843));
  OR2_X1    g418(.A1(G95), .A2(G2105), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n844), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT93), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G1991), .Z(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n738), .A2(G25), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n849), .B2(new_n852), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n840), .A2(new_n841), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT34), .ZN(new_n856));
  INV_X1    g431(.A(new_n609), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT81), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n610), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(G16), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT32), .B(G1981), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n779), .A2(G6), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n803), .A2(G22), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G303), .B2(new_n804), .ZN(new_n867));
  INV_X1    g442(.A(G1971), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n779), .B1(new_n581), .B2(new_n583), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n779), .A2(G23), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT33), .B(G1976), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT95), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n870), .B2(new_n872), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n867), .A2(new_n868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n864), .A2(new_n869), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n862), .B1(new_n860), .B2(new_n863), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n856), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n876), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n868), .B(new_n865), .C1(G166), .C2(new_n803), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n867), .A2(new_n868), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n881), .A2(new_n886), .A3(KEYINPUT34), .A4(new_n864), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n855), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT36), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI211_X1 g465(.A(KEYINPUT36), .B(new_n855), .C1(new_n880), .C2(new_n887), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n836), .B1(new_n890), .B2(new_n891), .ZN(G150));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n893));
  XNOR2_X1  g468(.A(G150), .B(new_n893), .ZN(G311));
  AOI22_X1  g469(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n511), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n554), .A2(G55), .A3(G543), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n554), .A2(G93), .A3(new_n509), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT102), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT102), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G860), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT37), .Z(new_n903));
  NOR2_X1   g478(.A1(new_n641), .A2(new_n654), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n656), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n556), .B(new_n896), .C1(new_n899), .C2(new_n900), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n906), .B(new_n909), .Z(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  INV_X1    g487(.A(G860), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n912), .B2(new_n914), .ZN(G145));
  XNOR2_X1  g490(.A(G162), .B(new_n481), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n668), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n848), .B(new_n675), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n751), .B(new_n761), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n489), .A2(G130), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT103), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n484), .A2(G142), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n468), .A2(G118), .ZN(new_n925));
  OAI21_X1  g500(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n814), .B(G164), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n927), .B(new_n928), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n919), .A2(new_n920), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n921), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n918), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n917), .A3(new_n931), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g514(.A1(new_n611), .A2(G166), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n858), .A2(G303), .A3(new_n859), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G288), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n626), .A2(new_n630), .A3(G288), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n940), .A2(new_n946), .A3(new_n947), .A4(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n909), .B(new_n659), .ZN(new_n954));
  NAND2_X1  g529(.A1(G299), .A2(new_n653), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n650), .A2(new_n641), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(G299), .A2(KEYINPUT104), .A3(new_n653), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(KEYINPUT41), .A3(new_n959), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT41), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n963), .A3(new_n957), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n954), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n953), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n953), .A3(new_n965), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n952), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n952), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n901), .A2(new_n657), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n971), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n901), .A2(new_n656), .ZN(new_n976));
  INV_X1    g551(.A(new_n908), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n545), .A2(G286), .A3(new_n546), .ZN(new_n978));
  AOI21_X1  g553(.A(G286), .B1(new_n545), .B2(new_n546), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NAND2_X1  g556(.A1(G171), .A2(G168), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n545), .A2(G286), .A3(new_n546), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n907), .A3(new_n908), .A4(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n909), .B(KEYINPUT106), .C1(new_n979), .C2(new_n978), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n962), .A2(new_n985), .A3(new_n964), .A4(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n958), .A2(new_n980), .A3(new_n959), .A4(new_n984), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n950), .A3(new_n949), .A4(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(new_n937), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n950), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT107), .B1(new_n949), .B2(new_n950), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n975), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n997));
  INV_X1    g572(.A(new_n950), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n940), .A2(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n960), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n985), .A2(new_n986), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n955), .A2(new_n957), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n980), .A2(new_n984), .B1(new_n1003), .B2(KEYINPUT41), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(KEYINPUT41), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1000), .A2(new_n992), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n989), .A2(new_n937), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT43), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n974), .B1(new_n996), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT108), .B1(new_n1011), .B2(KEYINPUT43), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n990), .A2(new_n995), .A3(new_n975), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(KEYINPUT44), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1010), .B1(new_n1012), .B2(new_n1015), .ZN(G397));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n499), .B2(new_n503), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n672), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1022));
  OAI21_X1  g597(.A(G40), .B1(new_n1022), .B2(new_n468), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n469), .A2(new_n471), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n479), .B2(G2105), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n472), .A2(KEYINPUT109), .A3(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n1017), .C1(new_n499), .C2(new_n503), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1020), .A2(new_n1025), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT111), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1020), .A4(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n868), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1031), .A2(new_n1037), .A3(new_n1034), .A4(new_n868), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1017), .C1(new_n499), .C2(new_n503), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1025), .A3(new_n1028), .A4(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1042), .A2(G2090), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1046));
  AND3_X1   g621(.A1(G303), .A2(G8), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(G303), .B2(G8), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(G8), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT115), .B(G1981), .Z(new_n1052));
  NAND4_X1  g627(.A1(new_n593), .A2(new_n601), .A3(new_n608), .A4(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n606), .A2(new_n592), .A3(new_n607), .A4(new_n589), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1018), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1032), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT49), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT116), .B(KEYINPUT49), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1056), .B(new_n1059), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n943), .A2(G1976), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1059), .A2(KEYINPUT114), .A3(KEYINPUT52), .A4(new_n1065), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n943), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1030), .A2(new_n786), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1032), .A2(new_n1074), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1077), .A2(new_n1057), .A3(G286), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1078), .A2(KEYINPUT63), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1049), .A2(new_n1051), .A3(new_n1072), .A4(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1039), .A2(new_n1084), .A3(new_n1025), .A4(new_n1028), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n745), .A3(new_n1041), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1057), .B1(new_n1035), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(new_n1050), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1051), .A2(new_n1072), .A3(new_n1088), .A4(new_n1078), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1080), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1064), .A2(new_n1094), .B1(new_n857), .B2(new_n1052), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1059), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1051), .A2(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1076), .B2(G286), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT123), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1073), .A2(new_n1075), .A3(new_n1100), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1103));
  OAI211_X1 g678(.A(G8), .B(new_n1102), .C1(new_n1103), .C2(G286), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1030), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1108), .A2(new_n1110), .B1(new_n1111), .B2(new_n1042), .ZN(new_n1112));
  AOI21_X1  g687(.A(G2078), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(KEYINPUT53), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1106), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1051), .A2(new_n1072), .A3(new_n1088), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1097), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1083), .A2(new_n1041), .A3(new_n1085), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1120), .A2(new_n1121), .B1(new_n1108), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n565), .B1(new_n647), .B2(new_n648), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(G299), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1119), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1085), .A2(new_n1041), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1084), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1121), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1108), .A2(new_n1122), .ZN(new_n1133));
  AND4_X1   g708(.A1(new_n1119), .A2(new_n1132), .A3(new_n1128), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1042), .A2(new_n782), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1032), .A2(new_n816), .A3(new_n1058), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n641), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1128), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT60), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1137), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n653), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(KEYINPUT122), .A3(new_n641), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1143), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1082), .B2(new_n1018), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1030), .B2(G1996), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n556), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT61), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT121), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1139), .A2(new_n1162), .A3(new_n1140), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1160), .B1(new_n1135), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1142), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1167));
  INV_X1    g742(.A(G2078), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1109), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1042), .A2(new_n1111), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1042), .A2(KEYINPUT124), .A3(new_n1111), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT53), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1023), .A2(new_n1024), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1020), .A2(new_n1029), .A3(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1173), .A2(new_n1174), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1170), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1173), .A2(new_n1174), .A3(new_n1179), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(G171), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1170), .A2(new_n1187), .A3(G301), .A4(new_n1112), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1112), .B(G301), .C1(new_n1113), .C2(KEYINPUT53), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT126), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1186), .A2(new_n1191), .A3(KEYINPUT54), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1103), .A2(G286), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1102), .A2(G8), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1193), .A2(new_n1194), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1170), .A2(new_n1180), .A3(G301), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1115), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT54), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1192), .A2(new_n1199), .A3(new_n1117), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1092), .B(new_n1118), .C1(new_n1166), .C2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n814), .B(new_n816), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT110), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n762), .ZN(new_n1204));
  INV_X1    g779(.A(G1996), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1082), .A2(new_n1020), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n848), .A2(new_n851), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n848), .A2(new_n851), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1207), .A2(new_n1205), .ZN(new_n1212));
  OAI211_X1 g787(.A(new_n1208), .B(new_n1211), .C1(new_n761), .C2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(G290), .B(G1986), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1201), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1212), .B(KEYINPUT46), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT47), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n626), .A2(new_n630), .A3(new_n838), .A4(new_n1207), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT48), .Z(new_n1222));
  OAI21_X1  g797(.A(new_n1220), .B1(new_n1213), .B2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1208), .B(new_n1210), .C1(new_n761), .C2(new_n1212), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1224), .B1(G2067), .B2(new_n814), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1223), .B1(new_n1207), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1216), .A2(new_n1226), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g802(.A1(new_n996), .A2(new_n1009), .ZN(new_n1229));
  INV_X1    g803(.A(G319), .ZN(new_n1230));
  NOR3_X1   g804(.A1(G401), .A2(new_n1230), .A3(G227), .ZN(new_n1231));
  OAI211_X1 g805(.A(new_n938), .B(new_n1231), .C1(new_n735), .C2(new_n736), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n1229), .A2(new_n1232), .ZN(G308));
  OAI21_X1  g807(.A(new_n1231), .B1(new_n735), .B2(new_n736), .ZN(new_n1234));
  AND3_X1   g808(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n1235));
  NOR2_X1   g809(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1236), .B1(new_n996), .B2(new_n1009), .ZN(G225));
endmodule


