//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332;
  XOR2_X1   g0000(.A(KEYINPUT65), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n205), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n203), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(G244), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n217), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n216), .B(new_n220), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  INV_X1    g0035(.A(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n223), .ZN(new_n239));
  XOR2_X1   g0039(.A(G226), .B(G232), .Z(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n211), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n202), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G223), .A2(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n213), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(G77), .C2(new_n253), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(new_n263), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n260), .B(new_n268), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n277), .A2(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n276), .A2(new_n284), .B1(new_n208), .B2(G20), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n276), .B2(new_n284), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n213), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(new_n271), .B2(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n275), .B(new_n295), .C1(new_n296), .C2(new_n274), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n268), .B1(new_n273), .B2(new_n228), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n253), .A2(G232), .A3(new_n254), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n307), .A2(new_n221), .A3(new_n254), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(G107), .B2(new_n307), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n298), .B(new_n300), .C1(new_n310), .C2(new_n270), .ZN(new_n311));
  INV_X1    g0111(.A(new_n288), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n315));
  INV_X1    g0115(.A(new_n277), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n282), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n292), .A2(G77), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G77), .B2(new_n290), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n310), .A2(new_n270), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n299), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n311), .B(new_n322), .C1(new_n324), .C2(G169), .ZN(new_n325));
  OAI211_X1 g0125(.A(G190), .B(new_n300), .C1(new_n310), .C2(new_n270), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n321), .B(new_n326), .C1(new_n324), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n274), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(G200), .B2(new_n274), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n297), .B(new_n329), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n279), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n282), .A2(G50), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n312), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT76), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT11), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT11), .ZN(new_n345));
  INV_X1    g0145(.A(new_n290), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT12), .B1(new_n346), .B2(new_n203), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n346), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n347), .B(new_n348), .C1(G68), .C2(new_n292), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT72), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n253), .A2(new_n355), .A3(G232), .A4(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(G226), .A3(new_n254), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT74), .A3(new_n259), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n363), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n354), .B2(new_n356), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n367), .B1(new_n369), .B2(new_n270), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n268), .B1(new_n273), .B2(new_n221), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT75), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n352), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  AOI211_X1 g0175(.A(KEYINPUT13), .B(new_n373), .C1(new_n366), .C2(new_n370), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n351), .B(G169), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT74), .B1(new_n365), .B2(new_n259), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n369), .A2(new_n367), .A3(new_n270), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n352), .A3(new_n374), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G179), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n351), .B1(new_n385), .B2(G169), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n350), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n350), .B1(new_n385), .B2(G200), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n330), .B2(new_n385), .ZN(new_n389));
  INV_X1    g0189(.A(new_n273), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(G232), .B1(new_n267), .B2(new_n264), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT77), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n305), .B2(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n278), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n306), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n269), .A2(G1698), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G223), .B2(G1698), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n392), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n259), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n391), .A2(new_n400), .A3(G190), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n327), .B1(new_n391), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n253), .B2(G20), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n305), .A2(G33), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT7), .B(new_n214), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n204), .A2(new_n206), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G20), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n282), .A2(G159), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n404), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n396), .A2(new_n405), .A3(new_n214), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n405), .B1(new_n396), .B2(new_n214), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n417), .A2(new_n418), .A3(new_n203), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n412), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT16), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n416), .B(new_n288), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n316), .A2(new_n290), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n292), .B2(new_n316), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n403), .A2(new_n422), .A3(KEYINPUT79), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n424), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n307), .B2(new_n214), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n405), .B(G20), .C1(new_n304), .C2(new_n306), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n420), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n312), .B1(new_n432), .B2(new_n404), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n396), .A2(new_n214), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n203), .B1(new_n434), .B2(KEYINPUT7), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n396), .A2(new_n405), .A3(new_n214), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT16), .A3(new_n420), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n428), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT79), .A3(KEYINPUT17), .A4(new_n403), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n427), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n399), .A2(new_n259), .ZN(new_n442));
  INV_X1    g0242(.A(G232), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n268), .B1(new_n273), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n391), .A2(new_n400), .A3(G179), .ZN(new_n446));
  AOI221_X4 g0246(.A(KEYINPUT18), .B1(new_n445), .B2(new_n446), .C1(new_n422), .C2(new_n424), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n416), .A2(new_n288), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n421), .B1(new_n436), .B2(new_n435), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n424), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n446), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT78), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n452), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT18), .B1(new_n439), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT78), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n448), .A3(new_n452), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n441), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n339), .A2(new_n387), .A3(new_n389), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G250), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n254), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT80), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(G33), .B2(G283), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n464), .A2(new_n307), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n394), .A2(new_n306), .A3(new_n395), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT4), .A2(G1698), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(G244), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n254), .A2(G244), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT4), .B1(new_n307), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n469), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT81), .B1(new_n475), .B2(new_n270), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n394), .A2(new_n395), .A3(G244), .A4(new_n306), .ZN(new_n477));
  INV_X1    g0277(.A(new_n471), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n469), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n259), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n271), .B(G45), .C1(new_n265), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G41), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n270), .B(G257), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(G41), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n271), .A4(G45), .ZN(new_n491));
  OAI21_X1  g0291(.A(G274), .B1(new_n258), .B2(new_n213), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT82), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n484), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n264), .A3(new_n495), .A4(new_n489), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n488), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n476), .A2(new_n483), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n502), .A2(new_n503), .A3(G107), .ZN(new_n504));
  XNOR2_X1  g0304(.A(G97), .B(G107), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n506), .A2(new_n214), .B1(new_n227), .B2(new_n283), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n406), .B2(new_n409), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n288), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n290), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n271), .A2(G33), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n213), .A2(new_n290), .A3(new_n287), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n493), .A2(new_n496), .B1(KEYINPUT83), .B2(new_n487), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n488), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n270), .B1(new_n479), .B2(new_n480), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(G190), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n488), .B(new_n516), .C1(new_n475), .C2(new_n270), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n296), .B1(new_n510), .B2(new_n514), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n476), .A2(new_n483), .A3(new_n298), .A4(new_n499), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n501), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n221), .A2(G1698), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n470), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n394), .A2(new_n395), .A3(new_n526), .A4(new_n306), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT85), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n477), .A2(new_n254), .B1(new_n278), .B2(new_n222), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n270), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n271), .B(G45), .C1(new_n534), .C2(G274), .ZN(new_n535));
  OAI211_X1 g0335(.A(KEYINPUT84), .B(G250), .C1(new_n266), .C2(G1), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n259), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n296), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n528), .B(new_n525), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n259), .B1(new_n539), .B2(new_n531), .ZN(new_n540));
  INV_X1    g0340(.A(new_n537), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n298), .A3(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n361), .A2(KEYINPUT19), .A3(new_n362), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n214), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n214), .A2(G68), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n396), .A2(new_n546), .B1(KEYINPUT19), .B2(new_n359), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n288), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n313), .A2(new_n346), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n513), .A2(new_n314), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n538), .A2(new_n542), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G200), .B1(new_n533), .B2(new_n537), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n540), .A2(G190), .A3(new_n541), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n513), .A2(G87), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n548), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(G20), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n470), .A2(KEYINPUT22), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n508), .A2(G20), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n508), .A3(G20), .ZN(new_n568));
  AOI22_X1  g0368(.A1(KEYINPUT90), .A2(new_n568), .B1(new_n279), .B2(G116), .ZN(new_n569));
  INV_X1    g0369(.A(new_n560), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n307), .A2(new_n570), .ZN(new_n571));
  OAI221_X1 g0371(.A(new_n569), .B1(KEYINPUT90), .B2(new_n568), .C1(new_n571), .C2(KEYINPUT22), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT24), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n569), .B1(KEYINPUT90), .B2(new_n568), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT22), .B1(new_n253), .B2(new_n560), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n563), .B(KEYINPUT89), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n561), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n312), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n508), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT91), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT25), .B1(new_n346), .B2(new_n508), .ZN(new_n583));
  XOR2_X1   g0383(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g0384(.A(new_n513), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n508), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n462), .A2(new_n254), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G257), .B2(new_n254), .ZN(new_n589));
  INV_X1    g0389(.A(G294), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n396), .A2(new_n589), .B1(new_n278), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n259), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n497), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n270), .B(G264), .C1(new_n484), .C2(new_n486), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT92), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT92), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n491), .A2(new_n596), .A3(G264), .A4(new_n270), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT93), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT93), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n593), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n592), .A3(new_n497), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n602), .A2(G200), .B1(G190), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n587), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n524), .A2(new_n558), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n290), .A2(G116), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n513), .B2(G116), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n214), .B1(new_n503), .B2(G33), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n465), .A2(KEYINPUT80), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n467), .A2(G33), .A3(G283), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n222), .A2(G20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n288), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(new_n278), .B2(G97), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n468), .B2(new_n466), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n287), .A2(new_n213), .B1(G20), .B2(new_n222), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n609), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n614), .B1(new_n613), .B2(new_n616), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n609), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n259), .B1(new_n494), .B2(new_n489), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n496), .A2(new_n493), .B1(new_n630), .B2(G270), .ZN(new_n631));
  OAI21_X1  g0431(.A(G303), .B1(new_n407), .B2(new_n408), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n236), .A2(G1698), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G257), .B2(G1698), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n396), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n259), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n296), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n607), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(G270), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n497), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n298), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n638), .A2(new_n639), .B1(new_n629), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n259), .A2(new_n591), .B1(new_n493), .B2(new_n496), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n595), .A2(new_n600), .A3(new_n597), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n600), .B1(new_n595), .B2(new_n597), .ZN(new_n646));
  OAI211_X1 g0446(.A(G179), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n603), .A2(G169), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n580), .B2(new_n586), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n641), .A2(G169), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n628), .B2(new_n623), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT21), .B1(new_n652), .B2(new_n607), .ZN(new_n653));
  INV_X1    g0453(.A(new_n629), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n641), .A2(G200), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n654), .B(new_n655), .C1(new_n330), .C2(new_n641), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n643), .A2(new_n650), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n461), .A2(new_n606), .A3(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n456), .A2(new_n458), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n375), .A2(new_n376), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT14), .B1(new_n661), .B2(new_n296), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n383), .A3(new_n377), .ZN(new_n663));
  INV_X1    g0463(.A(new_n325), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n350), .B1(new_n389), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n660), .B1(new_n665), .B2(new_n441), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n336), .A2(new_n338), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n297), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n552), .A2(new_n557), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n522), .A2(new_n523), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n629), .A2(new_n642), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n626), .A2(new_n627), .A3(new_n609), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n627), .B1(new_n626), .B2(new_n609), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n637), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(KEYINPUT87), .A3(new_n639), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n653), .A2(new_n650), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n587), .A2(new_n604), .B1(new_n501), .B2(new_n520), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n680), .B2(new_n670), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n672), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n552), .B(KEYINPUT94), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n668), .B1(new_n685), .B2(new_n461), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n643), .A2(new_n653), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n643), .A2(new_n653), .A3(new_n656), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n271), .A2(new_n214), .A3(G13), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n629), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g0495(.A(new_n687), .B(new_n688), .S(new_n695), .Z(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n694), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n587), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n605), .A3(new_n650), .ZN(new_n702));
  INV_X1    g0502(.A(new_n650), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n694), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n687), .A2(new_n699), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n694), .B(KEYINPUT96), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT97), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(KEYINPUT97), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n707), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n218), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n543), .A2(new_n222), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(G1), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n212), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n720), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  INV_X1    g0526(.A(new_n606), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n683), .B1(new_n727), .B2(new_n678), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n671), .B(KEYINPUT26), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n694), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  INV_X1    g0531(.A(new_n710), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n682), .B2(new_n684), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n733), .B2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n599), .A2(new_n601), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n642), .A2(new_n592), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n518), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n499), .A3(new_n540), .A4(new_n541), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n531), .B1(new_n527), .B2(new_n529), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n541), .B1(new_n741), .B2(new_n270), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n521), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n592), .B1(new_n645), .B2(new_n646), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n631), .A2(G179), .A3(new_n636), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(new_n746), .A3(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n641), .A2(new_n298), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n602), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT98), .A3(new_n500), .A4(new_n742), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT98), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n742), .A3(new_n298), .A4(new_n641), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n476), .A2(new_n483), .A3(new_n499), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n748), .A2(KEYINPUT99), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n751), .A3(new_n740), .A4(new_n747), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(new_n760), .A3(new_n694), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT31), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n657), .A2(new_n606), .A3(new_n732), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n748), .B1(new_n755), .B2(new_n754), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n732), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n763), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n734), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n726), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(G13), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G45), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n720), .A2(G1), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n697), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G330), .B2(new_n696), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n718), .A2(new_n307), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G355), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G116), .B2(new_n218), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n248), .A2(G45), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n470), .A2(new_n718), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n266), .B2(new_n212), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n782), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n262), .B1(new_n214), .B2(G169), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n777), .B1(new_n787), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT102), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n214), .A2(new_n298), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n798), .B1(new_n801), .B2(new_n330), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n800), .A2(KEYINPUT102), .A3(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G179), .A2(G200), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n214), .B1(new_n805), .B2(G190), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n203), .B1(new_n503), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT103), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n214), .A2(G190), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n805), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n800), .A2(new_n330), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n813), .C1(new_n815), .C2(new_n211), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n327), .A2(G179), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n809), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n508), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n214), .A2(new_n330), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n817), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(G87), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n298), .A2(G200), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n253), .C1(new_n227), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n820), .A2(new_n824), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT101), .Z(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n816), .B(new_n826), .C1(G58), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n808), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  INV_X1    g0632(.A(G326), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n307), .B1(new_n832), .B2(new_n821), .C1(new_n815), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n806), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(G294), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G283), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n818), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G322), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n827), .A2(new_n839), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n810), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n838), .B(new_n841), .C1(G329), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(KEYINPUT33), .B(G317), .Z(new_n844));
  OAI211_X1 g0644(.A(new_n836), .B(new_n843), .C1(new_n804), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n831), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n797), .B1(new_n846), .B2(new_n791), .ZN(new_n847));
  INV_X1    g0647(.A(new_n794), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n696), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n779), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  OAI21_X1  g0651(.A(new_n328), .B1(new_n321), .B2(new_n699), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n325), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n325), .A2(new_n694), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n733), .B(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n769), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n777), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(KEYINPUT105), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(KEYINPUT105), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n791), .A2(new_n792), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n776), .B1(new_n863), .B2(new_n227), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n253), .B1(new_n822), .B2(G107), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n865), .B1(new_n503), .B2(new_n806), .C1(new_n815), .C2(new_n832), .ZN(new_n866));
  INV_X1    g0666(.A(new_n827), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G294), .A2(new_n867), .B1(new_n842), .B2(G311), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n868), .B1(new_n559), .B2(new_n818), .C1(new_n222), .C2(new_n825), .ZN(new_n869));
  INV_X1    g0669(.A(new_n804), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n866), .B(new_n869), .C1(G283), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n825), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n829), .A2(G143), .B1(G159), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n870), .A2(G150), .B1(G137), .B2(new_n814), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT34), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n818), .A2(new_n203), .B1(new_n810), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n470), .B1(new_n202), .B2(new_n806), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n881), .B(new_n882), .C1(G50), .C2(new_n822), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n871), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n791), .ZN(new_n885));
  INV_X1    g0685(.A(new_n856), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n864), .B1(new_n884), .B2(new_n885), .C1(new_n886), .C2(new_n793), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n862), .A2(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n774), .A2(new_n271), .ZN(new_n889));
  INV_X1    g0689(.A(new_n441), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n447), .A2(new_n453), .A3(KEYINPUT78), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n457), .B1(new_n456), .B2(new_n458), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n450), .A2(new_n312), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n404), .B1(new_n419), .B2(new_n415), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n428), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n692), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT106), .B1(new_n460), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n439), .A2(new_n403), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n451), .A2(new_n452), .ZN(new_n904));
  INV_X1    g0704(.A(new_n692), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n451), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n903), .B1(new_n455), .B2(new_n897), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(new_n898), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n907), .B(KEYINPUT37), .Z(new_n915));
  AOI21_X1  g0715(.A(new_n906), .B1(new_n890), .B2(new_n660), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(KEYINPUT108), .A2(KEYINPUT39), .ZN(new_n919));
  AND2_X1   g0719(.A1(KEYINPUT108), .A2(KEYINPUT39), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n894), .B1(new_n893), .B2(new_n898), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n460), .A2(KEYINPUT106), .A3(new_n900), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n912), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n914), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n913), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT107), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(new_n925), .C2(new_n913), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n921), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n387), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n699), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n854), .B1(new_n733), .B2(new_n886), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n902), .B2(new_n912), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n914), .B(new_n911), .C1(new_n899), .C2(new_n901), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n350), .A2(new_n694), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n387), .A2(new_n389), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n663), .A2(new_n350), .A3(new_n694), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n934), .A2(new_n937), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n659), .B2(new_n692), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n461), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n731), .C1(new_n733), .C2(KEYINPUT29), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n668), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT109), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n945), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G330), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n757), .A2(new_n760), .A3(KEYINPUT31), .A4(new_n694), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n856), .B1(new_n939), .B2(new_n940), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n937), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT40), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n955), .A4(new_n956), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n461), .B1(new_n953), .B2(new_n954), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n961), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n889), .B1(new_n951), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n951), .B2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(new_n506), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(G116), .A3(new_n215), .A4(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT36), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n212), .A2(G77), .A3(new_n411), .ZN(new_n972));
  INV_X1    g0772(.A(new_n201), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n203), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(G1), .A3(new_n773), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n966), .A2(new_n971), .A3(new_n975), .ZN(G367));
  NAND2_X1  g0776(.A1(new_n732), .A2(new_n515), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n524), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n522), .A2(new_n523), .A3(new_n732), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n706), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT111), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n556), .A2(new_n699), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n683), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n669), .A2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n983), .B(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(new_n980), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n709), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT42), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n981), .A2(new_n703), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n732), .B1(new_n995), .B2(new_n670), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n991), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n990), .B(new_n998), .Z(new_n999));
  XOR2_X1   g0799(.A(new_n719), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT112), .B1(new_n716), .B2(new_n980), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n714), .A2(new_n1002), .A3(new_n715), .A4(new_n992), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(KEYINPUT44), .A3(new_n1003), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n992), .B1(new_n714), .B2(new_n715), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT45), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n707), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n705), .A2(new_n708), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n709), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n697), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1013), .A2(new_n771), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(KEYINPUT113), .A3(new_n706), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT113), .B1(new_n1017), .B2(new_n706), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1000), .B1(new_n1021), .B2(new_n771), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n775), .A2(G1), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n999), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n985), .A2(new_n848), .A3(new_n986), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n239), .A2(new_n785), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n795), .B1(new_n218), .B2(new_n313), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n777), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT114), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n814), .A2(G311), .B1(G107), .B2(new_n835), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT46), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n822), .A2(G116), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .C1(new_n804), .C2(new_n590), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n470), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(G317), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n825), .A2(new_n837), .B1(new_n810), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n818), .A2(new_n503), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1034), .B(new_n1038), .C1(new_n828), .C2(new_n832), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n806), .A2(new_n203), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n253), .B1(new_n818), .B2(new_n227), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G143), .C2(new_n814), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G58), .A2(new_n822), .B1(new_n842), .B2(G137), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n872), .A2(new_n973), .B1(new_n867), .B2(G150), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n804), .A2(new_n811), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1033), .A2(new_n1039), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT47), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n885), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1028), .A2(KEYINPUT114), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1029), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1025), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1024), .A2(new_n1054), .ZN(G387));
  NOR2_X1   g0855(.A1(new_n1014), .A2(new_n720), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n771), .B2(new_n1013), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n822), .A2(G294), .B1(new_n835), .B2(G283), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n814), .A2(G322), .B1(new_n872), .B2(G303), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n828), .B2(new_n1035), .C1(new_n804), .C2(new_n840), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT115), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT49), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n818), .A2(new_n222), .B1(new_n810), .B2(new_n833), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n470), .A3(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n825), .A2(new_n203), .B1(new_n810), .B2(new_n281), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G77), .B2(new_n822), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1037), .B1(G50), .B2(new_n867), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n814), .A2(G159), .B1(new_n314), .B2(new_n835), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1071), .A2(new_n470), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n316), .B2(new_n870), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n791), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n705), .A2(new_n794), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n780), .A2(new_n721), .B1(new_n508), .B2(new_n718), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n244), .A2(new_n266), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n316), .A2(new_n211), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT50), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n722), .B(new_n266), .C1(new_n203), .C2(new_n227), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n784), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n776), .B1(new_n1084), .B2(new_n795), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1076), .A2(new_n1077), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1057), .A2(new_n1058), .A3(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1017), .A2(new_n706), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1010), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1014), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1092), .B(new_n1014), .C1(new_n1088), .C2(new_n1010), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n719), .B(new_n1021), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1023), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n981), .A2(new_n848), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n795), .B1(new_n503), .B2(new_n218), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n785), .A2(new_n251), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n777), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n818), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G87), .A2(new_n1101), .B1(new_n842), .B2(G143), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n203), .B2(new_n821), .C1(new_n277), .C2(new_n825), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n806), .A2(new_n227), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n396), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n814), .A2(G150), .B1(new_n867), .B2(G159), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n201), .C2(new_n804), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n814), .A2(G317), .B1(new_n867), .B2(G311), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT52), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n870), .A2(G303), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n825), .A2(new_n590), .B1(new_n810), .B2(new_n839), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G283), .B2(new_n822), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n253), .B(new_n819), .C1(G116), .C2(new_n835), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1110), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1100), .B1(new_n1119), .B2(new_n791), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1096), .B1(new_n1097), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1094), .A2(new_n1121), .ZN(G390));
  NAND2_X1  g0922(.A1(new_n932), .A2(new_n699), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n934), .B2(new_n942), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n921), .B(new_n1124), .C1(new_n927), .C2(new_n930), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n854), .B1(new_n730), .B2(new_n853), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(new_n942), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1123), .A3(new_n918), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n768), .A2(new_n941), .A3(G330), .A4(new_n886), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n946), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n947), .A2(new_n668), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n768), .A2(G330), .A3(new_n886), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n942), .B1(new_n1131), .B2(new_n956), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(new_n1126), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n941), .B1(new_n1131), .B2(new_n886), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1136), .A2(new_n934), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT118), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n947), .A2(new_n668), .A3(new_n1140), .A4(new_n1132), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1134), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1128), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT39), .B1(new_n935), .B2(new_n936), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n928), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n926), .A2(KEYINPUT107), .A3(KEYINPUT39), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1143), .B1(new_n1148), .B2(new_n1124), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1131), .A2(new_n956), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1130), .B(new_n1142), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n956), .A3(new_n1131), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1130), .A4(new_n1142), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1130), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1142), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n720), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1154), .A2(new_n1023), .A3(new_n1130), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n863), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n777), .B1(new_n1163), .B2(new_n316), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n825), .A2(new_n1165), .B1(new_n806), .B2(new_n811), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n870), .B2(G137), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT120), .Z(new_n1168));
  NOR2_X1   g0968(.A1(new_n821), .A2(new_n281), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT53), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n814), .A2(G128), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n307), .B1(new_n842), .B2(G125), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1101), .A2(new_n973), .B1(new_n867), .B2(G132), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n870), .A2(G107), .B1(G97), .B2(new_n872), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT121), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n818), .A2(new_n203), .B1(new_n810), .B2(new_n590), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n867), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n307), .B1(new_n821), .B2(new_n559), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1104), .B(new_n1180), .C1(G283), .C2(new_n814), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1168), .A2(new_n1174), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1164), .B1(new_n1183), .B2(new_n791), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n931), .B2(new_n793), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1161), .A2(new_n1162), .A3(new_n1185), .ZN(G378));
  NAND2_X1  g0986(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G330), .B(new_n960), .C1(new_n958), .C2(KEYINPUT40), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n297), .B1(new_n336), .B2(new_n338), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n294), .A2(new_n905), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT55), .Z(new_n1192));
  XNOR2_X1  g0992(.A(new_n1190), .B(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1198));
  AND4_X1   g0998(.A1(new_n933), .A2(new_n1197), .A3(new_n944), .A4(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1197), .A2(new_n1198), .B1(new_n933), .B2(new_n944), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1188), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1188), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n719), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n777), .B1(new_n1163), .B2(new_n973), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n396), .B2(new_n265), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G107), .A2(new_n867), .B1(new_n1101), .B2(G58), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n837), .B2(new_n810), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1211), .A2(G41), .A3(new_n470), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n821), .A2(new_n227), .B1(new_n825), .B2(new_n313), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1040), .B(new_n1213), .C1(G116), .C2(new_n814), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(new_n503), .C2(new_n804), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(G128), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1218), .A2(new_n827), .B1(new_n821), .B2(new_n1165), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G137), .B2(new_n872), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n814), .A2(G125), .B1(G150), .B2(new_n835), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n804), .C2(new_n880), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1101), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n842), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1207), .B1(new_n1228), .B2(new_n791), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1195), .B2(new_n793), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT123), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1204), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n1023), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1206), .A2(new_n1233), .ZN(G375));
  INV_X1    g1034(.A(new_n1000), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1139), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1187), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1159), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n253), .B1(new_n1101), .B2(G77), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n313), .B2(new_n806), .C1(new_n815), .C2(new_n590), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G283), .A2(new_n867), .B1(new_n842), .B2(G303), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n503), .B2(new_n821), .C1(new_n508), .C2(new_n825), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G116), .C2(new_n870), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n829), .A2(G137), .B1(G132), .B2(new_n814), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n804), .B2(new_n1165), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G159), .A2(new_n822), .B1(new_n842), .B2(G128), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n202), .B2(new_n818), .C1(new_n281), .C2(new_n825), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n396), .B(new_n1248), .C1(G50), .C2(new_n835), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1243), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n777), .B1(G68), .B2(new_n1163), .C1(new_n1250), .C2(new_n885), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n942), .B2(new_n792), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1139), .B2(new_n1023), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1238), .A2(new_n1253), .ZN(G381));
  INV_X1    g1054(.A(new_n999), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT113), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1088), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1015), .B1(new_n1257), .B2(new_n1018), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1235), .B1(new_n1258), .B2(new_n770), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1259), .B2(new_n1095), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1260), .A2(G390), .A3(new_n1053), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(G375), .ZN(G407));
  NAND2_X1  g1065(.A1(new_n693), .A2(G213), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1262), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G407), .B(G213), .C1(G375), .C2(new_n1268), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1187), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1157), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1232), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n719), .B1(new_n1188), .B2(new_n1201), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1233), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT125), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1206), .A2(new_n1277), .A3(G378), .A4(new_n1233), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1095), .B1(new_n1188), .B2(new_n1000), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1232), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G378), .B1(new_n1281), .B2(new_n1230), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1159), .B(new_n719), .C1(new_n1285), .C2(new_n1237), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT60), .B1(new_n1187), .B2(new_n1236), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1253), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n862), .A3(new_n887), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1253), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1266), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1267), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1291), .B(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1282), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1267), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1293), .A2(new_n1294), .A3(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1024), .A2(new_n1054), .A3(new_n1094), .A4(new_n1121), .ZN(new_n1300));
  OAI21_X1  g1100(.A(G390), .B1(new_n1260), .B2(new_n1053), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(G393), .B(new_n850), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1300), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1297), .A2(new_n1267), .A3(new_n1291), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(KEYINPUT63), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1270), .B1(new_n1299), .B2(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1024), .A2(new_n1054), .B1(new_n1094), .B2(new_n1121), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1302), .B1(new_n1261), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1300), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1284), .A2(new_n1266), .A3(new_n1292), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1298), .A2(new_n1294), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(KEYINPUT126), .A4(new_n1293), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1309), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NOR4_X1   g1121(.A1(new_n1297), .A2(new_n1321), .A3(new_n1267), .A4(new_n1291), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1317), .B(KEYINPUT127), .C1(new_n1320), .C2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1313), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1327), .B2(new_n1317), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1319), .B1(new_n1324), .B2(new_n1328), .ZN(G405));
  AND2_X1   g1129(.A1(new_n1206), .A2(new_n1233), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1279), .B1(G378), .B2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1292), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1313), .ZN(G402));
endmodule


