//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  INV_X1    g004(.A(G50gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT14), .B(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n208), .A2(new_n214), .B1(KEYINPUT15), .B2(new_n202), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G8gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT91), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n226), .A2(new_n220), .A3(G8gat), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT17), .B1(new_n215), .B2(new_n216), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n230), .A3(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n235), .B(KEYINPUT13), .Z(new_n240));
  INV_X1    g039(.A(new_n236), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n217), .B1(new_n230), .B2(new_n231), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n238), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n234), .A2(new_n235), .A3(new_n236), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G169gat), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n243), .A3(new_n245), .A4(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G57gat), .B(G64gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT94), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260));
  NAND2_X1  g059(.A1(G71gat), .A2(G78gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(G71gat), .A2(G78gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT95), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  OR2_X1    g064(.A1(G57gat), .A2(G64gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G57gat), .A2(G64gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT94), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G71gat), .A2(G78gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G71gat), .A2(G78gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT95), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n262), .A2(new_n265), .A3(new_n268), .A4(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n261), .B(new_n263), .C1(new_n258), .C2(new_n260), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G231gat), .A2(G233gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G127gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G183gat), .B(G211gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n232), .B1(new_n275), .B2(new_n274), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT96), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n285), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n282), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT41), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT97), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n296), .B(KEYINPUT98), .Z(new_n297));
  XOR2_X1   g096(.A(G134gat), .B(G162gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G92gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n303));
  INV_X1    g102(.A(G85gat), .ZN(new_n304));
  OAI21_X1  g103(.A(G92gat), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT8), .ZN(new_n308));
  NAND2_X1  g107(.A1(G99gat), .A2(G106gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT99), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n310), .B2(new_n309), .ZN(new_n312));
  XNOR2_X1  g111(.A(G99gat), .B(G106gat), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n307), .B2(new_n312), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n219), .A2(new_n233), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G190gat), .B(G218gat), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n217), .A2(new_n316), .B1(KEYINPUT41), .B2(new_n294), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n318), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n300), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n299), .A3(new_n322), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n293), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n258), .A2(new_n259), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n261), .A2(new_n260), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n265), .A2(new_n268), .A3(new_n271), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n273), .ZN(new_n336));
  OAI22_X1  g135(.A1(new_n335), .A2(new_n336), .B1(new_n314), .B2(new_n315), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT10), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n307), .A2(new_n312), .ZN(new_n339));
  INV_X1    g138(.A(new_n313), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n341), .A2(new_n272), .A3(new_n273), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n316), .A2(KEYINPUT10), .A3(new_n273), .A4(new_n272), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n343), .ZN(new_n349));
  INV_X1    g148(.A(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT100), .ZN(new_n354));
  XNOR2_X1  g153(.A(G176gat), .B(G204gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(new_n351), .A3(new_n356), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n330), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT36), .ZN(new_n362));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT27), .B(G183gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT68), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n378), .A2(KEYINPUT26), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n378), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  INV_X1    g183(.A(G169gat), .ZN(new_n385));
  INV_X1    g184(.A(G176gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT23), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT65), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n377), .A2(new_n389), .A3(KEYINPUT23), .ZN(new_n390));
  INV_X1    g189(.A(new_n377), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT23), .B1(new_n385), .B2(new_n386), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n388), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  NAND4_X1  g194(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT64), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT25), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n392), .A2(new_n391), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT25), .A4(new_n387), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n384), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n387), .A2(KEYINPUT65), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n389), .B1(new_n377), .B2(KEYINPUT23), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(KEYINPUT66), .A3(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n383), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(G127gat), .A2(G134gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT69), .B(G127gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(G134gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(G113gat), .B2(G120gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G113gat), .ZN(new_n421));
  INV_X1    g220(.A(G120gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n415), .ZN(new_n425));
  NAND2_X1  g224(.A1(G127gat), .A2(G134gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n419), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT70), .B(G113gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G120gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT71), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n414), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n417), .A2(new_n423), .B1(new_n427), .B2(new_n429), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n383), .B(new_n435), .C1(new_n406), .C2(new_n413), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n364), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(G15gat), .B(G43gat), .Z(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n446));
  INV_X1    g245(.A(new_n435), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n401), .A2(new_n405), .A3(new_n384), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT66), .B1(new_n412), .B2(new_n404), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n414), .B2(new_n432), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n451), .B2(new_n364), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n414), .A2(new_n432), .ZN(new_n453));
  NAND2_X1  g252(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n363), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n443), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n437), .B(KEYINPUT32), .C1(new_n439), .C2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n444), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n438), .A2(new_n440), .A3(new_n443), .ZN(new_n460));
  INV_X1    g259(.A(new_n458), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT73), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT73), .B1(new_n452), .B2(new_n455), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n464), .B2(KEYINPUT74), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  OAI221_X1 g265(.A(new_n466), .B1(new_n462), .B2(new_n463), .C1(new_n460), .C2(new_n461), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n362), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT31), .B(G50gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G211gat), .B(G218gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT22), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT75), .B(G211gat), .Z(new_n472));
  INV_X1    g271(.A(G218gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G197gat), .B(G204gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n470), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G141gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G148gat), .ZN(new_n482));
  INV_X1    g281(.A(G148gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G141gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G155gat), .B(G162gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT2), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(G155gat), .A2(G162gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(G155gat), .A2(G162gat), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT77), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G162gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n287), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n487), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n492), .A2(new_n496), .B1(new_n485), .B2(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT3), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n483), .A2(G141gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n481), .A2(G148gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n488), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT77), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n495), .B1(new_n494), .B2(new_n487), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n499), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G228gat), .ZN(new_n512));
  INV_X1    g311(.A(G233gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n503), .B(new_n498), .C1(new_n504), .C2(new_n505), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n497), .A2(new_n498), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n478), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n474), .A2(new_n523), .A3(new_n470), .A4(new_n475), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(new_n509), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n521), .B1(new_n526), .B2(new_n500), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n478), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n509), .B1(new_n529), .B2(new_n476), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n521), .B1(new_n530), .B2(new_n500), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n515), .B1(new_n532), .B2(new_n511), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n469), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n479), .B1(new_n509), .B2(new_n508), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n514), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n469), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(new_n516), .C2(new_n527), .ZN(new_n538));
  XNOR2_X1  g337(.A(G78gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G22gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n534), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n534), .B2(new_n538), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G1gat), .B(G29gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G85gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT5), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n431), .B1(new_n519), .B2(new_n520), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n499), .A2(new_n507), .A3(new_n434), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G225gat), .A2(G233gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n499), .A2(new_n507), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT79), .B1(new_n558), .B2(KEYINPUT3), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n508), .A2(new_n431), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n500), .B1(new_n499), .B2(new_n507), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n555), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n552), .B2(KEYINPUT4), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT4), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n499), .A2(new_n568), .A3(new_n507), .A4(new_n434), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT81), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n521), .A2(new_n571), .A3(new_n568), .A4(new_n434), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n565), .A3(KEYINPUT4), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n567), .A2(new_n570), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n557), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n431), .B(new_n508), .C1(new_n562), .C2(KEYINPUT79), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n550), .B(new_n554), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n552), .A2(KEYINPUT4), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n569), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n568), .A4(new_n434), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n549), .B1(new_n575), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n572), .A2(new_n570), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n552), .A2(new_n565), .A3(KEYINPUT4), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n586), .A2(new_n566), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n554), .B1(new_n576), .B2(new_n577), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n556), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n581), .A2(new_n582), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n564), .A2(new_n591), .A3(new_n550), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n548), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT6), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(KEYINPUT6), .B(new_n549), .C1(new_n575), .C2(new_n584), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G8gat), .B(G36gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G64gat), .B(G92gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(G226gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n513), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n446), .B(new_n602), .C1(new_n401), .C2(new_n405), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(KEYINPUT29), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n480), .B(new_n603), .C1(new_n414), .C2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n446), .B1(new_n401), .B2(new_n405), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n414), .A2(new_n602), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n608), .B2(new_n480), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT76), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT76), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n611), .C1(new_n608), .C2(new_n480), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n600), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n606), .B(new_n600), .C1(new_n608), .C2(new_n480), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT30), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n604), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n618));
  INV_X1    g417(.A(new_n602), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n479), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n621), .A2(KEYINPUT30), .A3(new_n606), .A4(new_n600), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n543), .B1(new_n597), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n459), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n452), .A2(new_n455), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n460), .B2(new_n461), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n626), .A2(new_n362), .A3(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n468), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT87), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n581), .B(new_n582), .C1(new_n576), .C2(new_n577), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n555), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n548), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT39), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT85), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n555), .B2(new_n633), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n632), .B1(new_n636), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n585), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n633), .A2(new_n555), .ZN(new_n646));
  INV_X1    g445(.A(new_n641), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT85), .B1(new_n637), .B2(KEYINPUT39), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(KEYINPUT40), .A3(new_n548), .A4(new_n635), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n613), .B2(new_n623), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n543), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n614), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n606), .B(new_n655), .C1(new_n608), .C2(new_n480), .ZN(new_n656));
  INV_X1    g455(.A(new_n600), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n603), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n618), .B2(new_n604), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n660), .B2(new_n479), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n620), .A2(new_n480), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT38), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n654), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n595), .A2(new_n664), .A3(new_n596), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n610), .A2(new_n612), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT37), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n665), .A2(KEYINPUT86), .B1(KEYINPUT38), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT86), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n595), .A2(new_n664), .A3(new_n670), .A4(new_n596), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n631), .B(new_n653), .C1(new_n669), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(KEYINPUT86), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(KEYINPUT38), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n653), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT87), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n630), .B1(new_n672), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n465), .A2(new_n467), .A3(new_n543), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n597), .A2(new_n624), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT35), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n541), .A2(new_n542), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n626), .A2(new_n628), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n597), .A4(new_n624), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n257), .B(new_n361), .C1(new_n678), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n597), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(G1gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1324gat));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  INV_X1    g492(.A(new_n624), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT102), .Z(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(G8gat), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n695), .A2(new_n693), .A3(new_n697), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(G1325gat));
  AOI21_X1  g500(.A(G15gat), .B1(new_n688), .B2(new_n685), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n468), .A2(new_n629), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT103), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n688), .B2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n682), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  AOI21_X1  g508(.A(new_n328), .B1(new_n678), .B2(new_n687), .ZN(new_n710));
  INV_X1    g509(.A(new_n293), .ZN(new_n711));
  INV_X1    g510(.A(new_n360), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n257), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n212), .A3(new_n689), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(new_n687), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n678), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n630), .B(KEYINPUT104), .C1(new_n672), .C2(new_n677), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n328), .A2(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n722), .A2(new_n724), .B1(new_n725), .B2(new_n710), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n713), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n597), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n717), .A2(new_n728), .ZN(G1328gat));
  AOI21_X1  g528(.A(G36gat), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n694), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n727), .B2(new_n624), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  NAND2_X1  g534(.A1(new_n703), .A2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n685), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n727), .A2(new_n736), .B1(G43gat), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g539(.A(new_n206), .B1(new_n714), .B2(new_n543), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n682), .A2(G50gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n727), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g543(.A1(new_n330), .A2(new_n257), .A3(new_n712), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n689), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g547(.A1(new_n722), .A2(new_n624), .A3(new_n745), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n703), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n737), .A2(G71gat), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n754), .A2(G71gat), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n746), .A2(new_n682), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n711), .A2(new_n256), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n712), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n726), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n597), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n675), .A2(new_n676), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n631), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n675), .A2(KEYINPUT87), .A3(new_n676), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT104), .B1(new_n768), .B2(new_n630), .ZN(new_n769));
  INV_X1    g568(.A(new_n721), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n687), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n760), .A2(new_n329), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n722), .B2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n689), .A2(new_n304), .A3(new_n712), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT106), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n764), .B1(new_n778), .B2(new_n780), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n624), .A2(new_n360), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n771), .B2(new_n773), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n722), .A2(new_n775), .A3(new_n772), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n301), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n624), .A2(new_n301), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n720), .A2(new_n721), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n724), .B1(new_n792), .B2(new_n687), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n710), .A2(new_n725), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n762), .B(new_n791), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n783), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n785), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(G92gat), .B1(new_n777), .B2(new_n786), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n784), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(G1337gat));
  INV_X1    g601(.A(new_n703), .ZN(new_n803));
  OAI21_X1  g602(.A(G99gat), .B1(new_n763), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n737), .A2(G99gat), .A3(new_n360), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT108), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n778), .B2(new_n806), .ZN(G1338gat));
  OAI211_X1 g606(.A(new_n682), .B(new_n762), .C1(new_n793), .C2(new_n794), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n543), .A2(G106gat), .A3(new_n360), .ZN(new_n810));
  OAI211_X1 g609(.A(KEYINPUT109), .B(new_n810), .C1(new_n787), .C2(new_n788), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT109), .B1(new_n777), .B2(new_n810), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n726), .A2(new_n816), .A3(new_n682), .A4(new_n762), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n817), .A3(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n777), .B2(new_n810), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n346), .B2(new_n347), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT54), .B(new_n350), .C1(new_n344), .C2(new_n345), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(KEYINPUT111), .A3(new_n356), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n346), .A2(new_n823), .A3(new_n347), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n357), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n826), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n359), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT111), .B1(new_n827), .B2(new_n356), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n829), .A3(new_n357), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n824), .A2(new_n825), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT112), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n828), .B2(new_n831), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n822), .ZN(new_n841));
  INV_X1    g640(.A(new_n359), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n836), .B2(new_n826), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n256), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n241), .A2(new_n242), .A3(new_n240), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n251), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n712), .A2(new_n255), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n329), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n255), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n255), .B2(new_n849), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n328), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n839), .A3(new_n845), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n293), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n330), .A2(new_n257), .A3(new_n360), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n597), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n679), .A2(new_n694), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n257), .A2(new_n428), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n859), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT114), .B1(new_n865), .B2(new_n543), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(new_n682), .C1(new_n858), .C2(new_n859), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n689), .A2(new_n869), .A3(new_n624), .A4(new_n685), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n256), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n864), .B1(new_n872), .B2(new_n421), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n862), .B2(new_n712), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n360), .A2(new_n422), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n870), .B2(new_n875), .ZN(G1341gat));
  INV_X1    g675(.A(new_n416), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n870), .B2(new_n711), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n862), .A2(new_n877), .A3(new_n711), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n862), .A2(new_n881), .A3(new_n329), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n881), .B1(new_n870), .B2(new_n329), .ZN(new_n887));
  OR3_X1    g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G1343gat));
  XNOR2_X1  g687(.A(new_n850), .B(KEYINPUT116), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n841), .A2(new_n843), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n257), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n328), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n856), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n293), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n859), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n893), .B2(new_n293), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n682), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT57), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n543), .B1(new_n858), .B2(new_n859), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n703), .A2(new_n597), .A3(new_n694), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n257), .ZN(new_n905));
  AND4_X1   g704(.A1(new_n682), .A2(new_n860), .A3(new_n624), .A4(new_n803), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n481), .A3(new_n256), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT58), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n905), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n906), .A2(new_n483), .A3(new_n712), .ZN(new_n913));
  INV_X1    g712(.A(new_n904), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT59), .B(new_n483), .C1(new_n914), .C2(new_n712), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n900), .A2(new_n901), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n890), .A2(KEYINPUT118), .A3(new_n328), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n853), .A2(new_n854), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT118), .B1(new_n890), .B2(new_n328), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n711), .B1(new_n892), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n859), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n901), .B(new_n682), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n712), .A3(new_n903), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n913), .B1(new_n915), .B2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n904), .B2(new_n293), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n906), .A2(new_n287), .A3(new_n711), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  AOI21_X1  g730(.A(G162gat), .B1(new_n906), .B2(new_n329), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n328), .A2(new_n493), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n914), .B2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n689), .A2(new_n624), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n679), .B(new_n936), .C1(new_n858), .C2(new_n859), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n385), .A3(new_n256), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT119), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n936), .A2(new_n737), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n869), .A2(new_n256), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n942), .B2(new_n385), .ZN(G1348gat));
  NAND2_X1  g742(.A1(new_n869), .A2(new_n940), .ZN(new_n944));
  OAI21_X1  g743(.A(G176gat), .B1(new_n944), .B2(new_n360), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n937), .A2(new_n386), .A3(new_n712), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  NOR2_X1   g746(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n948));
  OAI21_X1  g747(.A(G183gat), .B1(new_n944), .B2(new_n293), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n373), .A3(new_n711), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1350gat));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n329), .B(new_n940), .C1(new_n866), .C2(new_n868), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n956), .A2(G190gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT121), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n963));
  XNOR2_X1  g762(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n937), .A2(new_n370), .A3(new_n329), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n960), .A2(new_n965), .A3(KEYINPUT123), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n703), .A2(new_n936), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n925), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n256), .A2(G197gat), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n900), .A2(new_n972), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(new_n256), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n973), .A2(new_n974), .B1(G197gat), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(G1352gat));
  OAI21_X1  g777(.A(G204gat), .B1(new_n973), .B2(new_n360), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(G204gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n975), .A2(new_n981), .A3(new_n712), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n982), .A2(new_n984), .A3(KEYINPUT62), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n982), .B2(KEYINPUT62), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n985), .A2(new_n986), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n979), .A4(new_n983), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(new_n991), .ZN(G1353gat));
  OAI21_X1  g791(.A(KEYINPUT126), .B1(new_n973), .B2(new_n293), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n925), .A2(new_n994), .A3(new_n711), .A4(new_n972), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n993), .A2(G211gat), .A3(new_n995), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT63), .ZN(new_n998));
  XNOR2_X1  g797(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n993), .A2(G211gat), .A3(new_n995), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n975), .A2(new_n472), .A3(new_n711), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n973), .B2(new_n328), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n975), .A2(new_n473), .A3(new_n329), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1355gat));
endmodule


