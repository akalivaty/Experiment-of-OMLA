

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(G2104), .A2(n518), .ZN(n873) );
  AND2_X2 U547 ( .A1(n518), .A2(G2104), .ZN(n869) );
  OR2_X1 U548 ( .A1(n514), .A2(n647), .ZN(n637) );
  XNOR2_X1 U549 ( .A(n669), .B(n668), .ZN(n671) );
  INV_X1 U550 ( .A(KEYINPUT64), .ZN(n668) );
  INV_X1 U551 ( .A(KEYINPUT33), .ZN(n670) );
  OR2_X1 U552 ( .A1(n596), .A2(n513), .ZN(n597) );
  NOR2_X1 U553 ( .A1(n616), .A2(n615), .ZN(n625) );
  NOR2_X1 U554 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U555 ( .A1(n662), .A2(n661), .ZN(n680) );
  NAND2_X1 U556 ( .A1(n671), .A2(n670), .ZN(n676) );
  NAND2_X1 U557 ( .A1(n709), .A2(n593), .ZN(n653) );
  AND2_X1 U558 ( .A1(n653), .A2(G1341), .ZN(n513) );
  OR2_X1 U559 ( .A1(n648), .A2(n636), .ZN(n514) );
  INV_X1 U560 ( .A(G8), .ZN(n636) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n630) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n642) );
  INV_X1 U563 ( .A(n708), .ZN(n593) );
  NAND2_X1 U564 ( .A1(G8), .A2(n653), .ZN(n685) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  NOR2_X1 U566 ( .A1(n558), .A2(G651), .ZN(n780) );
  NOR2_X1 U567 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U568 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U569 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U570 ( .A1(G126), .A2(n873), .ZN(n516) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U572 ( .A1(G114), .A2(n874), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U574 ( .A(n517), .B(KEYINPUT83), .ZN(n521) );
  NAND2_X1 U575 ( .A1(G102), .A2(n869), .ZN(n519) );
  XNOR2_X1 U576 ( .A(n519), .B(KEYINPUT84), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n521), .A2(n520), .ZN(n525) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n522), .Z(n870) );
  NAND2_X1 U579 ( .A1(G138), .A2(n870), .ZN(n523) );
  XNOR2_X1 U580 ( .A(KEYINPUT85), .B(n523), .ZN(n524) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n558) );
  NAND2_X1 U582 ( .A1(n780), .A2(G52), .ZN(n530) );
  INV_X1 U583 ( .A(G651), .ZN(n531) );
  NOR2_X1 U584 ( .A1(G543), .A2(n531), .ZN(n527) );
  XNOR2_X1 U585 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n526) );
  XNOR2_X1 U586 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U587 ( .A(KEYINPUT67), .B(n528), .ZN(n781) );
  NAND2_X1 U588 ( .A1(G64), .A2(n781), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n784) );
  NAND2_X1 U591 ( .A1(G90), .A2(n784), .ZN(n533) );
  NOR2_X1 U592 ( .A1(n558), .A2(n531), .ZN(n785) );
  NAND2_X1 U593 ( .A1(G77), .A2(n785), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n534), .Z(n535) );
  NOR2_X1 U596 ( .A1(n536), .A2(n535), .ZN(G171) );
  NAND2_X1 U597 ( .A1(n784), .A2(G89), .ZN(n537) );
  XNOR2_X1 U598 ( .A(n537), .B(KEYINPUT4), .ZN(n539) );
  NAND2_X1 U599 ( .A1(G76), .A2(n785), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n540), .B(KEYINPUT5), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n780), .A2(G51), .ZN(n542) );
  NAND2_X1 U603 ( .A1(G63), .A2(n781), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(n780), .A2(G50), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G62), .A2(n781), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G88), .A2(n784), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G75), .A2(n785), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT77), .B(n551), .Z(n552) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(G166) );
  XOR2_X1 U617 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U618 ( .A1(G49), .A2(n780), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G74), .A2(G651), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT76), .B(n556), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n781), .A2(n557), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n558), .A2(G87), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(G288) );
  NAND2_X1 U625 ( .A1(n784), .A2(G86), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G61), .A2(n781), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n785), .A2(G73), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT2), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n780), .A2(G48), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(G305) );
  NAND2_X1 U633 ( .A1(G85), .A2(n784), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G72), .A2(n785), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n780), .A2(G47), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G60), .A2(n781), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  OR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(G290) );
  NOR2_X1 U640 ( .A1(G164), .A2(G1384), .ZN(n709) );
  NAND2_X1 U641 ( .A1(G101), .A2(n869), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT66), .ZN(n576) );
  INV_X1 U643 ( .A(KEYINPUT23), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G125), .A2(n873), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G137), .A2(n870), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G113), .A2(n874), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U650 ( .A(KEYINPUT65), .B(n583), .Z(n743) );
  NAND2_X1 U651 ( .A1(n743), .A2(G40), .ZN(n708) );
  NOR2_X1 U652 ( .A1(G1966), .A2(n685), .ZN(n647) );
  NAND2_X1 U653 ( .A1(n781), .A2(G56), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n584), .Z(n590) );
  NAND2_X1 U655 ( .A1(n784), .A2(G81), .ZN(n585) );
  XNOR2_X1 U656 ( .A(n585), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G68), .A2(n785), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n588), .Z(n589) );
  NOR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n780), .A2(G43), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n991) );
  AND2_X1 U663 ( .A1(n709), .A2(n593), .ZN(n594) );
  AND2_X1 U664 ( .A1(n594), .A2(G1996), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n595), .B(KEYINPUT26), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n991), .A2(n597), .ZN(n609) );
  NAND2_X1 U667 ( .A1(G79), .A2(n785), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G54), .A2(n780), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n604) );
  NAND2_X1 U670 ( .A1(n784), .A2(G92), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G66), .A2(n781), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(KEYINPUT72), .B(n602), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT15), .ZN(n987) );
  NAND2_X1 U676 ( .A1(G1348), .A2(n653), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G2067), .A2(n594), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n610) );
  NOR2_X1 U679 ( .A1(n987), .A2(n610), .ZN(n608) );
  OR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n987), .A2(n610), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n624) );
  NAND2_X1 U683 ( .A1(G1956), .A2(n653), .ZN(n613) );
  XNOR2_X1 U684 ( .A(KEYINPUT93), .B(n613), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n594), .A2(G2072), .ZN(n614) );
  XNOR2_X1 U686 ( .A(KEYINPUT27), .B(n614), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n780), .A2(G53), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G65), .A2(n781), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G91), .A2(n784), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G78), .A2(n785), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n980) );
  NAND2_X1 U694 ( .A1(n625), .A2(n980), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n629) );
  NOR2_X1 U696 ( .A1(n625), .A2(n980), .ZN(n627) );
  XOR2_X1 U697 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(n635) );
  OR2_X1 U701 ( .A1(n594), .A2(G1961), .ZN(n633) );
  XNOR2_X1 U702 ( .A(G2078), .B(KEYINPUT25), .ZN(n942) );
  NAND2_X1 U703 ( .A1(n594), .A2(n942), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n639) );
  NAND2_X1 U705 ( .A1(n639), .A2(G171), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n645) );
  NOR2_X1 U707 ( .A1(G2084), .A2(n653), .ZN(n648) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT30), .ZN(n638) );
  NOR2_X1 U709 ( .A1(G168), .A2(n638), .ZN(n641) );
  NOR2_X1 U710 ( .A1(G171), .A2(n639), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n652) );
  XNOR2_X1 U713 ( .A(KEYINPUT95), .B(n652), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U715 ( .A1(G8), .A2(n648), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n662) );
  AND2_X1 U717 ( .A1(G286), .A2(G8), .ZN(n651) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n659) );
  NOR2_X1 U719 ( .A1(G1971), .A2(n685), .ZN(n655) );
  NOR2_X1 U720 ( .A1(G2090), .A2(n653), .ZN(n654) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U722 ( .A1(n656), .A2(G303), .ZN(n657) );
  OR2_X1 U723 ( .A1(n636), .A2(n657), .ZN(n658) );
  AND2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U725 ( .A(KEYINPUT32), .B(n660), .ZN(n661) );
  NOR2_X1 U726 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NOR2_X1 U727 ( .A1(G303), .A2(G1971), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n979), .A2(n663), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n680), .A2(n664), .ZN(n667) );
  NAND2_X1 U730 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U731 ( .A(n981), .ZN(n665) );
  NOR2_X1 U732 ( .A1(n665), .A2(n685), .ZN(n666) );
  AND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n979), .A2(KEYINPUT33), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n672), .A2(n685), .ZN(n674) );
  XOR2_X1 U736 ( .A(G1981), .B(G305), .Z(n996) );
  INV_X1 U737 ( .A(n996), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT96), .ZN(n689) );
  NOR2_X1 U741 ( .A1(G2090), .A2(G303), .ZN(n678) );
  NAND2_X1 U742 ( .A1(G8), .A2(n678), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U744 ( .A(KEYINPUT97), .B(n681), .Z(n682) );
  AND2_X1 U745 ( .A1(n682), .A2(n685), .ZN(n687) );
  NOR2_X1 U746 ( .A1(G1981), .A2(G305), .ZN(n683) );
  XOR2_X1 U747 ( .A(n683), .B(KEYINPUT24), .Z(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  AND2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n724) );
  XOR2_X1 U751 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n691) );
  NAND2_X1 U752 ( .A1(G105), .A2(n869), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(n695) );
  NAND2_X1 U754 ( .A1(G129), .A2(n873), .ZN(n693) );
  NAND2_X1 U755 ( .A1(G141), .A2(n870), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n874), .A2(G117), .ZN(n696) );
  NAND2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n865) );
  NAND2_X1 U760 ( .A1(G1996), .A2(n865), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT91), .ZN(n707) );
  INV_X1 U762 ( .A(G1991), .ZN(n936) );
  NAND2_X1 U763 ( .A1(G107), .A2(n874), .ZN(n700) );
  NAND2_X1 U764 ( .A1(G95), .A2(n869), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U766 ( .A1(G119), .A2(n873), .ZN(n702) );
  NAND2_X1 U767 ( .A1(G131), .A2(n870), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U770 ( .A(n705), .B(KEYINPUT89), .Z(n880) );
  NOR2_X1 U771 ( .A1(n936), .A2(n880), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n917) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n738) );
  XOR2_X1 U774 ( .A(n738), .B(KEYINPUT92), .Z(n710) );
  NOR2_X1 U775 ( .A1(n917), .A2(n710), .ZN(n730) );
  INV_X1 U776 ( .A(n730), .ZN(n722) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n736) );
  NAND2_X1 U778 ( .A1(n870), .A2(G140), .ZN(n711) );
  XOR2_X1 U779 ( .A(KEYINPUT87), .B(n711), .Z(n713) );
  NAND2_X1 U780 ( .A1(n869), .A2(G104), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U782 ( .A(KEYINPUT34), .B(n714), .ZN(n720) );
  NAND2_X1 U783 ( .A1(G128), .A2(n873), .ZN(n716) );
  NAND2_X1 U784 ( .A1(G116), .A2(n874), .ZN(n715) );
  NAND2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U786 ( .A(KEYINPUT35), .B(n717), .Z(n718) );
  XNOR2_X1 U787 ( .A(KEYINPUT88), .B(n718), .ZN(n719) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U789 ( .A(KEYINPUT36), .B(n721), .ZN(n887) );
  NOR2_X1 U790 ( .A1(n736), .A2(n887), .ZN(n926) );
  NAND2_X1 U791 ( .A1(n738), .A2(n926), .ZN(n734) );
  NAND2_X1 U792 ( .A1(n722), .A2(n734), .ZN(n723) );
  NOR2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U794 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U795 ( .A1(n993), .A2(n738), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n741) );
  XOR2_X1 U797 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n733) );
  NOR2_X1 U798 ( .A1(G1996), .A2(n865), .ZN(n919) );
  AND2_X1 U799 ( .A1(n880), .A2(n936), .ZN(n727) );
  XNOR2_X1 U800 ( .A(n727), .B(KEYINPUT98), .ZN(n915) );
  NOR2_X1 U801 ( .A1(G1986), .A2(G290), .ZN(n728) );
  NOR2_X1 U802 ( .A1(n915), .A2(n728), .ZN(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U804 ( .A1(n919), .A2(n731), .ZN(n732) );
  XNOR2_X1 U805 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n736), .A2(n887), .ZN(n923) );
  NAND2_X1 U808 ( .A1(n737), .A2(n923), .ZN(n739) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U811 ( .A(n742), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U812 ( .A(n743), .Z(G160) );
  XNOR2_X1 U813 ( .A(G2451), .B(G2435), .ZN(n753) );
  XOR2_X1 U814 ( .A(G2446), .B(KEYINPUT101), .Z(n745) );
  XNOR2_X1 U815 ( .A(G2454), .B(G2430), .ZN(n744) );
  XNOR2_X1 U816 ( .A(n745), .B(n744), .ZN(n749) );
  XOR2_X1 U817 ( .A(KEYINPUT100), .B(G2427), .Z(n747) );
  XNOR2_X1 U818 ( .A(G1341), .B(G1348), .ZN(n746) );
  XNOR2_X1 U819 ( .A(n747), .B(n746), .ZN(n748) );
  XOR2_X1 U820 ( .A(n749), .B(n748), .Z(n751) );
  XNOR2_X1 U821 ( .A(G2443), .B(G2438), .ZN(n750) );
  XNOR2_X1 U822 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U823 ( .A(n753), .B(n752), .ZN(n754) );
  AND2_X1 U824 ( .A1(n754), .A2(G14), .ZN(G401) );
  AND2_X1 U825 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U826 ( .A(G57), .ZN(G237) );
  NAND2_X1 U827 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U828 ( .A(n755), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U829 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n757) );
  XNOR2_X1 U830 ( .A(G223), .B(KEYINPUT69), .ZN(n821) );
  NAND2_X1 U831 ( .A1(G567), .A2(n821), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n757), .B(n756), .ZN(G234) );
  INV_X1 U833 ( .A(G860), .ZN(n764) );
  OR2_X1 U834 ( .A1(n991), .A2(n764), .ZN(G153) );
  XNOR2_X1 U835 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U836 ( .A1(G868), .A2(G301), .ZN(n759) );
  INV_X1 U837 ( .A(G868), .ZN(n761) );
  NAND2_X1 U838 ( .A1(n987), .A2(n761), .ZN(n758) );
  NAND2_X1 U839 ( .A1(n759), .A2(n758), .ZN(G284) );
  INV_X1 U840 ( .A(n980), .ZN(G299) );
  NOR2_X1 U841 ( .A1(G868), .A2(G299), .ZN(n760) );
  XOR2_X1 U842 ( .A(KEYINPUT73), .B(n760), .Z(n763) );
  NOR2_X1 U843 ( .A1(G286), .A2(n761), .ZN(n762) );
  NOR2_X1 U844 ( .A1(n763), .A2(n762), .ZN(G297) );
  NAND2_X1 U845 ( .A1(n764), .A2(G559), .ZN(n765) );
  INV_X1 U846 ( .A(n987), .ZN(n790) );
  NAND2_X1 U847 ( .A1(n765), .A2(n790), .ZN(n766) );
  XNOR2_X1 U848 ( .A(n766), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U849 ( .A1(G868), .A2(n991), .ZN(n769) );
  NAND2_X1 U850 ( .A1(n790), .A2(G868), .ZN(n767) );
  NOR2_X1 U851 ( .A1(G559), .A2(n767), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(G282) );
  NAND2_X1 U853 ( .A1(n873), .A2(G123), .ZN(n770) );
  XNOR2_X1 U854 ( .A(n770), .B(KEYINPUT18), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G135), .A2(n870), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U857 ( .A(KEYINPUT74), .B(n773), .ZN(n777) );
  NAND2_X1 U858 ( .A1(G111), .A2(n874), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G99), .A2(n869), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n911) );
  XNOR2_X1 U862 ( .A(n911), .B(G2096), .ZN(n779) );
  INV_X1 U863 ( .A(G2100), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(G156) );
  NAND2_X1 U865 ( .A1(n780), .A2(G55), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G67), .A2(n781), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G93), .A2(n784), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G80), .A2(n785), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U871 ( .A1(n789), .A2(n788), .ZN(n799) );
  NAND2_X1 U872 ( .A1(G559), .A2(n790), .ZN(n791) );
  XNOR2_X1 U873 ( .A(n791), .B(n991), .ZN(n802) );
  NOR2_X1 U874 ( .A1(G860), .A2(n802), .ZN(n792) );
  XOR2_X1 U875 ( .A(KEYINPUT75), .B(n792), .Z(n793) );
  XNOR2_X1 U876 ( .A(n799), .B(n793), .ZN(G145) );
  NOR2_X1 U877 ( .A1(G868), .A2(n799), .ZN(n794) );
  XNOR2_X1 U878 ( .A(n794), .B(KEYINPUT79), .ZN(n805) );
  XNOR2_X1 U879 ( .A(n980), .B(KEYINPUT78), .ZN(n795) );
  XNOR2_X1 U880 ( .A(n795), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U881 ( .A(G166), .B(G305), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n796), .B(G288), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n798), .B(n797), .ZN(n801) );
  XNOR2_X1 U884 ( .A(G290), .B(n799), .ZN(n800) );
  XNOR2_X1 U885 ( .A(n801), .B(n800), .ZN(n890) );
  XNOR2_X1 U886 ( .A(n890), .B(n802), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G868), .A2(n803), .ZN(n804) );
  NAND2_X1 U888 ( .A1(n805), .A2(n804), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n806) );
  XOR2_X1 U890 ( .A(KEYINPUT20), .B(n806), .Z(n807) );
  NAND2_X1 U891 ( .A1(G2090), .A2(n807), .ZN(n808) );
  XNOR2_X1 U892 ( .A(KEYINPUT21), .B(n808), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n809), .A2(G2072), .ZN(n810) );
  XNOR2_X1 U894 ( .A(KEYINPUT80), .B(n810), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U896 ( .A1(G69), .A2(G120), .ZN(n811) );
  NOR2_X1 U897 ( .A1(G237), .A2(n811), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G108), .A2(n812), .ZN(n826) );
  NAND2_X1 U899 ( .A1(n826), .A2(G567), .ZN(n819) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n814) );
  NAND2_X1 U901 ( .A1(G132), .A2(G82), .ZN(n813) );
  XNOR2_X1 U902 ( .A(n814), .B(n813), .ZN(n815) );
  NOR2_X1 U903 ( .A1(n815), .A2(G218), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G96), .A2(n816), .ZN(n825) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n825), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT82), .B(n817), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n819), .A2(n818), .ZN(n827) );
  NAND2_X1 U908 ( .A1(G483), .A2(G661), .ZN(n820) );
  NOR2_X1 U909 ( .A1(n827), .A2(n820), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U917 ( .A(G132), .ZN(G219) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G82), .ZN(G220) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n827), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2100), .B(KEYINPUT103), .Z(n829) );
  XNOR2_X1 U926 ( .A(G2678), .B(KEYINPUT102), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2090), .Z(n831) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT42), .B(G2096), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U934 ( .A(G2084), .B(G2078), .Z(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1961), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n840), .B(G2474), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1981), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1966), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G112), .A2(n874), .ZN(n848) );
  NAND2_X1 U947 ( .A1(G100), .A2(n869), .ZN(n847) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n856) );
  XOR2_X1 U949 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n850) );
  NAND2_X1 U950 ( .A1(G124), .A2(n873), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT104), .B(n851), .ZN(n854) );
  NAND2_X1 U953 ( .A1(G136), .A2(n870), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n852), .B(KEYINPUT106), .ZN(n853) );
  NAND2_X1 U955 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U957 ( .A1(G130), .A2(n873), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G118), .A2(n874), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G106), .A2(n869), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G142), .A2(n870), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n911), .B(n864), .ZN(n886) );
  XNOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT107), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(G160), .B(n868), .ZN(n884) );
  NAND2_X1 U970 ( .A1(G103), .A2(n869), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G127), .A2(n873), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n906) );
  XOR2_X1 U978 ( .A(n906), .B(G162), .Z(n882) );
  XNOR2_X1 U979 ( .A(G164), .B(n880), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U983 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U984 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U985 ( .A(G286), .B(n890), .ZN(n893) );
  XOR2_X1 U986 ( .A(G171), .B(KEYINPUT108), .Z(n891) );
  XNOR2_X1 U987 ( .A(n991), .B(n891), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(n987), .B(n894), .Z(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT109), .B(n896), .Z(G397) );
  NOR2_X1 U992 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n899), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(KEYINPUT112), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G401), .A2(n903), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n904), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  INV_X1 U1002 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1003 ( .A(G164), .B(G2078), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT113), .ZN(n908) );
  XOR2_X1 U1005 ( .A(G2072), .B(n906), .Z(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT50), .B(n909), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G2084), .B(G160), .Z(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n922) );
  XOR2_X1 U1013 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n920), .B(KEYINPUT51), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1019 ( .A(KEYINPUT52), .B(n927), .ZN(n929) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1022 ( .A1(n930), .A2(G29), .ZN(n1013) );
  XOR2_X1 U1023 ( .A(G2090), .B(G35), .Z(n933) );
  XOR2_X1 U1024 ( .A(G34), .B(KEYINPUT54), .Z(n931) );
  XNOR2_X1 U1025 ( .A(G2084), .B(n931), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n947) );
  XNOR2_X1 U1027 ( .A(G1996), .B(G32), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(G33), .B(G2072), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(G25), .B(n936), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(G28), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G26), .B(G2067), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n944) );
  XOR2_X1 U1035 ( .A(G27), .B(n942), .Z(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n945), .B(KEYINPUT53), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(n948), .Z(n949) );
  XNOR2_X1 U1040 ( .A(KEYINPUT114), .B(n949), .ZN(n950) );
  NOR2_X1 U1041 ( .A1(G29), .A2(n950), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT115), .B(n951), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n952), .A2(G11), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(n953), .B(KEYINPUT116), .ZN(n1011) );
  XNOR2_X1 U1045 ( .A(G21), .B(G1966), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n954), .B(KEYINPUT123), .ZN(n974) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(G1341), .B(G19), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G6), .B(G1981), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT121), .B(n957), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT122), .B(n960), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G1348), .B(KEYINPUT59), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(G4), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n964), .B(KEYINPUT60), .ZN(n972) );
  XNOR2_X1 U1058 ( .A(G1986), .B(G24), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G1971), .B(G22), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1061 ( .A(G1976), .B(KEYINPUT124), .Z(n967) );
  XNOR2_X1 U1062 ( .A(G23), .B(n967), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G5), .B(G1961), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT61), .B(n977), .Z(n978) );
  NOR2_X1 U1070 ( .A1(G16), .A2(n978), .ZN(n1008) );
  XNOR2_X1 U1071 ( .A(KEYINPUT56), .B(G16), .ZN(n1005) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT119), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1956), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G303), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G1348), .B(n987), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT118), .B(n988), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n1003) );
  XNOR2_X1 U1081 ( .A(G171), .B(G1961), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n991), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT57), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n999), .B(KEYINPUT117), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(KEYINPUT120), .B(n1006), .Z(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(n1009), .B(KEYINPUT125), .ZN(n1010) );
  NOR2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(KEYINPUT62), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1015), .ZN(G150) );
  INV_X1 U1099 ( .A(G150), .ZN(G311) );
endmodule

