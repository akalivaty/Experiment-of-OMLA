//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1077, new_n1078;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(new_n466), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n466), .A2(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(G136), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  INV_X1    g059(.A(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT3), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G126), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n466), .A2(new_n491), .A3(G126), .A4(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n465), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT70), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  AOI211_X1 g074(.A(new_n499), .B(new_n496), .C1(new_n490), .C2(new_n492), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n466), .A2(G138), .A3(new_n465), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n484), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NOR4_X1   g083(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT71), .A4(new_n506), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(G543), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT72), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n530), .B2(new_n521), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT73), .Z(new_n532));
  INV_X1    g107(.A(new_n524), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(G51), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT74), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n521), .A2(new_n540), .B1(new_n541), .B2(new_n524), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n518), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(new_n549), .B1(G43), .B2(new_n533), .ZN(new_n550));
  INV_X1    g125(.A(new_n521), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  XNOR2_X1  g135(.A(KEYINPUT76), .B(G65), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n516), .A2(new_n561), .B1(G78), .B2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT77), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(G91), .B2(new_n551), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n533), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n551), .A2(G87), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT78), .Z(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n533), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n516), .A2(KEYINPUT79), .A3(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n515), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G86), .B2(new_n551), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n533), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n518), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n521), .A2(new_n586), .B1(new_n587), .B2(new_n524), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n551), .A2(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n518), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n533), .A2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G321));
  XNOR2_X1  g175(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n553), .A2(new_n602), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n598), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n474), .A2(G123), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT81), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n479), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT82), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n479), .A2(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XOR2_X1   g201(.A(G2443), .B(G2446), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n630), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT17), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(KEYINPUT18), .B2(new_n642), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n648), .B(new_n651), .Z(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n654), .B2(new_n658), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G1991), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  OAI21_X1  g250(.A(KEYINPUT88), .B1(G16), .B2(G23), .ZN(new_n676));
  OR3_X1    g251(.A1(KEYINPUT88), .A2(G16), .A3(G23), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n677), .C1(G288), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT33), .B(G1976), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(KEYINPUT89), .B1(new_n683), .B2(G16), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n683), .A2(KEYINPUT89), .A3(G16), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(G166), .C2(new_n678), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G1971), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n681), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(G1971), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n678), .A2(G6), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n678), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT32), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT90), .Z(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n479), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n474), .A2(G119), .ZN(new_n700));
  NOR2_X1   g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G25), .B(new_n703), .S(G29), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT35), .B(G1991), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT87), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n678), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n589), .B2(new_n678), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(new_n667), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n697), .A2(new_n698), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2090), .ZN(new_n718));
  INV_X1    g293(.A(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT92), .B1(new_n719), .B2(G16), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n719), .A2(KEYINPUT92), .A3(G16), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n720), .B(new_n721), .C1(new_n554), .C2(new_n678), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1341), .Z(new_n723));
  INV_X1    g298(.A(G299), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT23), .B1(new_n724), .B2(new_n678), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n678), .A2(G20), .ZN(new_n726));
  MUX2_X1   g301(.A(KEYINPUT23), .B(new_n725), .S(new_n726), .Z(new_n727));
  OAI21_X1  g302(.A(new_n723), .B1(new_n727), .B2(G1956), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G1956), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n678), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n678), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1966), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n678), .A2(G4), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n599), .B2(new_n678), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2072), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n714), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n479), .A2(G139), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT95), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n743), .C1(new_n465), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(G29), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n618), .A2(G29), .B1(new_n737), .B2(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(G141), .A2(new_n479), .B1(new_n474), .B2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n756), .A2(new_n714), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G160), .B2(new_n714), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(G2084), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT30), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n759), .B2(G2084), .ZN(new_n764));
  INV_X1    g339(.A(new_n746), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2072), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n736), .A2(new_n747), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G171), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G5), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n772));
  INV_X1    g347(.A(G26), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n776));
  INV_X1    g351(.A(G104), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n465), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n474), .A2(G128), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n479), .A2(G140), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(G29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n772), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n769), .A2(new_n770), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(G2067), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n771), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n732), .A2(new_n767), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n714), .A2(KEYINPUT96), .A3(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n714), .ZN(new_n791));
  AOI21_X1  g366(.A(KEYINPUT96), .B1(new_n714), .B2(G27), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT97), .B(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT31), .B(G11), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n729), .A2(new_n789), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n713), .A2(new_n718), .A3(new_n797), .ZN(G311));
  INV_X1    g373(.A(G311), .ZN(G150));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n521), .A2(new_n800), .B1(new_n801), .B2(new_n524), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n516), .A2(G67), .ZN(new_n803));
  NAND2_X1  g378(.A1(G80), .A2(G543), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n518), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G860), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT37), .Z(new_n809));
  OAI21_X1  g384(.A(new_n553), .B1(KEYINPUT98), .B2(new_n806), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n810), .B(new_n811), .Z(new_n812));
  NOR2_X1   g387(.A1(new_n598), .A2(new_n606), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n812), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n809), .B1(new_n816), .B2(G860), .ZN(G145));
  OR2_X1    g392(.A1(new_n506), .A2(KEYINPUT99), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n496), .B1(new_n490), .B2(new_n492), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n506), .A2(KEYINPUT99), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n782), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n752), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n745), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n479), .A2(G142), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n474), .A2(G130), .ZN(new_n827));
  NOR2_X1   g402(.A1(G106), .A2(G2105), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n703), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT100), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n621), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n825), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(KEYINPUT101), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n834), .B(KEYINPUT102), .C1(new_n835), .C2(new_n824), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n618), .B(G162), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G160), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g417(.A1(new_n807), .A2(new_n602), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n812), .B(new_n609), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n724), .B(new_n598), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT41), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(new_n844), .ZN(new_n848));
  XNOR2_X1  g423(.A(G166), .B(new_n589), .ZN(new_n849));
  XNOR2_X1  g424(.A(G288), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G305), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(KEYINPUT103), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n848), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n843), .B1(new_n856), .B2(new_n602), .ZN(G331));
  XNOR2_X1  g432(.A(G331), .B(KEYINPUT104), .ZN(G295));
  XNOR2_X1  g433(.A(G168), .B(G171), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(new_n812), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n812), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n846), .ZN(new_n863));
  MUX2_X1   g438(.A(new_n862), .B(new_n860), .S(KEYINPUT105), .Z(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(new_n845), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n865), .B2(new_n854), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n864), .A2(new_n846), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n845), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n854), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n866), .B1(new_n854), .B2(new_n865), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n871), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT106), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n867), .A2(new_n870), .ZN(new_n875));
  MUX2_X1   g450(.A(new_n875), .B(new_n872), .S(KEYINPUT43), .Z(new_n876));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(G397));
  INV_X1    g454(.A(G2067), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n782), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G1996), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n752), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n703), .A2(new_n705), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n884), .A2(new_n885), .B1(G2067), .B2(new_n782), .ZN(new_n886));
  INV_X1    g461(.A(G1384), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n821), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n889));
  NAND2_X1  g464(.A1(G160), .A2(G40), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n881), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n895), .B2(new_n752), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(KEYINPUT46), .A3(new_n882), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n892), .B2(G1996), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT47), .Z(new_n901));
  INV_X1    g476(.A(new_n884), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n885), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n703), .B2(new_n705), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n892), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT125), .Z(new_n906));
  NOR2_X1   g481(.A1(G290), .A2(G1986), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n893), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT48), .ZN(new_n909));
  AOI211_X1 g484(.A(new_n894), .B(new_n901), .C1(new_n906), .C2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n510), .A2(KEYINPUT113), .A3(KEYINPUT45), .A4(new_n887), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n890), .B1(new_n888), .B2(new_n889), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n493), .A2(new_n497), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n499), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n819), .A2(KEYINPUT70), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n507), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT71), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n484), .A3(new_n507), .A4(new_n915), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(KEYINPUT45), .A3(new_n887), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(new_n912), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1966), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT114), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n887), .A3(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n888), .A2(KEYINPUT50), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n891), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(G2084), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n931), .A3(new_n923), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT119), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT119), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n925), .A2(new_n935), .A3(new_n930), .A4(new_n932), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(G8), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n937), .A2(KEYINPUT120), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT120), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(new_n939), .A3(G8), .A4(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(G8), .ZN(new_n941));
  NOR2_X1   g516(.A1(G168), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT51), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT121), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT121), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(KEYINPUT51), .C1(new_n938), .C2(new_n944), .ZN(new_n948));
  AOI211_X1 g523(.A(KEYINPUT51), .B(new_n942), .C1(new_n933), .C2(G8), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT122), .Z(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n934), .A2(new_n942), .A3(new_n936), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n821), .A2(KEYINPUT45), .A3(new_n887), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT107), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n890), .B1(new_n926), .B2(new_n889), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(G1971), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n958), .B2(G1971), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n960), .B(new_n962), .C1(G2090), .C2(new_n929), .ZN(new_n963));
  NAND2_X1  g538(.A1(G303), .A2(G8), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT55), .Z(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(G8), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n888), .A2(new_n890), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n941), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(G288), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n968), .B(KEYINPUT109), .C1(new_n969), .C2(G288), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n972), .B(new_n973), .Z(new_n974));
  AOI21_X1  g549(.A(KEYINPUT110), .B1(new_n580), .B2(G651), .ZN(new_n975));
  INV_X1    g550(.A(G1981), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(G305), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(KEYINPUT111), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n968), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n974), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n888), .A2(KEYINPUT50), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n891), .C1(new_n926), .C2(KEYINPUT50), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G2090), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n959), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n965), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n966), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2078), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n958), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT123), .B(G1961), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n929), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(KEYINPUT53), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n922), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n993), .A2(G171), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n951), .A2(new_n1001), .A3(new_n952), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n954), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G301), .B(KEYINPUT54), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n956), .A2(KEYINPUT53), .A3(new_n994), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1006), .B2(new_n912), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n992), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT56), .B(G2072), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n956), .A2(new_n957), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1956), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n987), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT57), .B1(new_n564), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n724), .B(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT61), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n929), .A2(new_n735), .B1(new_n880), .B2(new_n967), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(new_n598), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n598), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1021), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1023), .A3(new_n599), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n958), .A2(new_n1031), .A3(new_n882), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT58), .B(G1341), .Z(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n888), .B2(new_n890), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n956), .A2(new_n957), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT116), .B1(new_n1035), .B2(G1996), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n554), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(KEYINPUT117), .B2(KEYINPUT59), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1040), .B(new_n1038), .C1(new_n1039), .C2(KEYINPUT59), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1019), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1025), .A2(new_n1020), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1009), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n951), .B2(new_n952), .ZN(new_n1047));
  INV_X1    g622(.A(new_n966), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(new_n985), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n691), .A2(new_n976), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT112), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n984), .A2(new_n969), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(G288), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n968), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n933), .A2(G8), .A3(G168), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT63), .B1(new_n993), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n966), .A2(new_n985), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n965), .B1(new_n963), .B2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NOR4_X1   g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1055), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1054), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1047), .A2(new_n1049), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1003), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n904), .B1(new_n667), .B2(new_n589), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n893), .B1(new_n1065), .B2(new_n907), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT124), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1066), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1068), .B(new_n1069), .C1(new_n1003), .C2(new_n1063), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n910), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT126), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT126), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n910), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g650(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1077));
  XOR2_X1   g651(.A(new_n1077), .B(KEYINPUT127), .Z(new_n1078));
  NAND3_X1  g652(.A1(new_n876), .A2(new_n841), .A3(new_n1078), .ZN(G225));
  INV_X1    g653(.A(G225), .ZN(G308));
endmodule


