//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(new_n449), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n468), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT71), .B1(new_n467), .B2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND4_X1  g055(.A1(new_n475), .A2(new_n472), .A3(G2105), .A4(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(G136), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n474), .A2(G114), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(new_n490), .A3(KEYINPUT72), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n494), .A2(new_n496), .B1(new_n481), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n475), .A2(new_n472), .A3(new_n468), .A4(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n466), .A2(new_n468), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n498), .A2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .A3(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n508), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n513), .A2(G651), .B1(G50), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(new_n510), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT74), .B(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n524), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n511), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n515), .B1(new_n540), .B2(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n521), .A2(G90), .A3(new_n522), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n545), .A2(KEYINPUT77), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT77), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n515), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n521), .A2(G81), .A3(new_n522), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n521), .A2(G43), .A3(G543), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT78), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT78), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AND3_X1   g138(.A1(new_n521), .A2(G91), .A3(new_n522), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n509), .A2(new_n565), .A3(new_n510), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n565), .B1(new_n509), .B2(new_n510), .ZN(new_n568));
  OAI21_X1  g143(.A(G65), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n564), .B1(new_n571), .B2(G651), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT80), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n522), .A2(KEYINPUT79), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n566), .ZN(new_n578));
  INV_X1    g153(.A(new_n570), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n564), .ZN(new_n581));
  AND4_X1   g156(.A1(KEYINPUT80), .A2(new_n574), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n575), .A2(new_n582), .ZN(G299));
  NAND2_X1  g158(.A1(new_n524), .A2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n519), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n511), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n524), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n524), .A2(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n519), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT81), .B(G47), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n594), .B1(new_n515), .B2(new_n595), .C1(new_n596), .C2(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(new_n521), .A2(G92), .A3(new_n522), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n577), .B2(new_n566), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT82), .Z(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n519), .A2(G54), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n601), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G284));
  XOR2_X1   g186(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  XNOR2_X1  g190(.A(G280), .B(KEYINPUT84), .ZN(G297));
  INV_X1    g191(.A(G860), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n608), .B1(G559), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT85), .ZN(G148));
  NAND2_X1  g194(.A1(new_n557), .A2(new_n609), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n608), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g198(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n467), .A2(new_n465), .A3(G2105), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n629));
  OAI22_X1  g204(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(G2100), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n628), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n474), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI22_X1  g211(.A1(new_n481), .A2(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n487), .B2(G135), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT88), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT89), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(new_n681), .B(new_n680), .S(new_n673), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1986), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n687), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n687), .B2(new_n691), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(KEYINPUT101), .A2(KEYINPUT26), .ZN(new_n702));
  NAND2_X1  g277(.A1(KEYINPUT101), .A2(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n477), .A2(G105), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G129), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n487), .A2(G141), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT102), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n705), .B(new_n706), .C1(new_n708), .C2(new_n481), .ZN(new_n714));
  INV_X1    g289(.A(G141), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n486), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(G32), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  INV_X1    g300(.A(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n726), .B2(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(KEYINPUT24), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n479), .B2(new_n720), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n720), .A2(G33), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n487), .A2(G139), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n466), .A2(new_n468), .ZN(new_n735));
  INV_X1    g310(.A(G127), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n733), .B1(G2105), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT100), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(KEYINPUT100), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n730), .B1(new_n744), .B2(new_n720), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n724), .B1(new_n725), .B2(new_n729), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT103), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n752), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT104), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT29), .B(G2090), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n720), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n720), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n761), .B1(G2078), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G2078), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G171), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G5), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n759), .A2(new_n760), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n729), .A2(new_n725), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT31), .B(G11), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n777), .A2(KEYINPUT105), .B1(KEYINPUT30), .B2(new_n775), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n638), .B2(G29), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n772), .A2(new_n773), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n770), .A2(new_n771), .A3(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n766), .B(new_n783), .C1(new_n722), .C2(new_n723), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n752), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n614), .B2(new_n752), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n752), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n558), .B2(new_n752), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT98), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n608), .B2(new_n752), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1348), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n720), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT28), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n800));
  INV_X1    g375(.A(G128), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n481), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n487), .B2(G140), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(new_n720), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n792), .A2(new_n796), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT99), .Z(new_n808));
  NAND3_X1  g383(.A1(new_n751), .A2(new_n789), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n720), .A2(G25), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(KEYINPUT92), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(KEYINPUT92), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  INV_X1    g391(.A(G119), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n481), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n487), .A2(G131), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g396(.A(new_n811), .B(new_n812), .C1(new_n821), .C2(G29), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n752), .A2(G24), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G290), .B2(G16), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(new_n688), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n688), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n822), .A2(new_n823), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n591), .A2(G16), .A3(new_n592), .ZN(new_n831));
  OR2_X1    g406(.A1(G6), .A2(G16), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT32), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G1981), .ZN(new_n838));
  INV_X1    g413(.A(G1981), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(G303), .A2(G16), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n752), .A2(G22), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT94), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G1971), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(G1971), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n752), .A2(G23), .ZN(new_n852));
  INV_X1    g427(.A(G288), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n752), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT33), .B(G1976), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n841), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n829), .B(new_n830), .C1(new_n857), .C2(KEYINPUT34), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT95), .B1(new_n857), .B2(KEYINPUT34), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(KEYINPUT95), .A3(KEYINPUT34), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT97), .Z(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n862), .B2(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n809), .B1(new_n869), .B2(new_n871), .ZN(G311));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n871), .ZN(new_n873));
  INV_X1    g448(.A(new_n809), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(G150));
  AOI22_X1  g450(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n876), .A2(new_n515), .B1(new_n523), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n519), .A2(G55), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(new_n617), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  INV_X1    g457(.A(new_n608), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G559), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n878), .A2(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n557), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n554), .A2(new_n553), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT78), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n554), .A2(new_n553), .A3(KEYINPUT78), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n552), .A3(new_n880), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n885), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT106), .Z(new_n898));
  OAI21_X1  g473(.A(new_n617), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n882), .B1(new_n898), .B2(new_n899), .ZN(G145));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n498), .B2(new_n504), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n498), .A2(new_n504), .A3(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT102), .B1(new_n710), .B2(new_n711), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n714), .A2(new_n716), .A3(new_n713), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n902), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n712), .B(new_n717), .C1(new_n908), .C2(new_n903), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n907), .A2(new_n909), .A3(new_n803), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n803), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT108), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n740), .B1(new_n912), .B2(new_n741), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n909), .ZN(new_n914));
  INV_X1    g489(.A(new_n803), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n907), .A2(new_n909), .A3(new_n803), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n743), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G130), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n474), .A2(G118), .ZN(new_n922));
  OAI21_X1  g497(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n481), .A2(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n487), .B2(G142), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n820), .B(new_n925), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n627), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n913), .A2(new_n920), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n926), .B(new_n626), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n916), .A2(new_n918), .A3(new_n917), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n739), .B1(new_n930), .B2(KEYINPUT100), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n931), .B2(new_n919), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(KEYINPUT109), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n638), .B(new_n479), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(G162), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n936), .B(new_n929), .C1(new_n931), .C2(new_n919), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT110), .B(G37), .Z(new_n939));
  XOR2_X1   g514(.A(new_n935), .B(KEYINPUT111), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n930), .A2(KEYINPUT100), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n919), .B1(new_n941), .B2(new_n740), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(new_n927), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n932), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n938), .A2(KEYINPUT40), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT40), .B1(new_n938), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(G395));
  OAI21_X1  g522(.A(KEYINPUT114), .B1(new_n880), .B2(G868), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n608), .B1(new_n575), .B2(new_n582), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n574), .A2(new_n580), .A3(new_n581), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT80), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n572), .A2(KEYINPUT80), .A3(new_n574), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n883), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(KEYINPUT112), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  NAND3_X1  g531(.A1(G299), .A2(new_n956), .A3(new_n883), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(KEYINPUT41), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(new_n959), .A3(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n894), .B(new_n621), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(G305), .B(G303), .Z(new_n964));
  XNOR2_X1  g539(.A(G290), .B(new_n853), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n966), .A2(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n957), .B2(new_n955), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n963), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n962), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n958), .B2(new_n960), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n970), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n968), .A2(new_n969), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n609), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n948), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n971), .B1(new_n963), .B2(new_n973), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n976), .A2(new_n970), .A3(new_n972), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n984), .A2(new_n987), .A3(G868), .A4(new_n982), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n983), .A2(new_n988), .ZN(G295));
  NOR2_X1   g564(.A1(new_n983), .A2(new_n988), .ZN(G331));
  NAND3_X1  g565(.A1(new_n887), .A2(G301), .A3(new_n893), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(G301), .B1(new_n887), .B2(new_n893), .ZN(new_n993));
  OAI21_X1  g568(.A(G286), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n894), .A2(G171), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G168), .A3(new_n991), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n994), .A2(new_n996), .B1(new_n955), .B2(new_n957), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n996), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n961), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n966), .A2(new_n967), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n998), .B1(new_n958), .B2(new_n960), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1004), .B2(new_n997), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n949), .A2(new_n954), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n999), .A2(KEYINPUT41), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n994), .A2(KEYINPUT41), .A3(new_n996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n955), .A2(new_n957), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n939), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1012), .A2(new_n1005), .A3(KEYINPUT43), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT44), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1005), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1015), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1019), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g595(.A(G1996), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n718), .B(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n803), .B(G2067), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n820), .B(new_n823), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n498), .B2(new_n504), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n470), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1032), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G290), .B(new_n688), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1031), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT45), .B(new_n1027), .C1(new_n498), .C2(new_n504), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1041), .A2(new_n1030), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1031), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(new_n1043), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1044), .A2(new_n1046), .A3(G1971), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1031), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(new_n1027), .C1(new_n498), .C2(new_n504), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1048), .A2(KEYINPUT117), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(new_n1040), .C1(new_n1047), .C2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n853), .A2(G1976), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n591), .A2(new_n839), .A3(new_n592), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n839), .B1(new_n591), .B2(new_n592), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1065), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(new_n1060), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1060), .A2(new_n1061), .A3(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1063), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1057), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1030), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT116), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1045), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1052), .B1(new_n1080), .B2(G1971), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1040), .B1(new_n1081), .B2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n769), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1045), .A2(KEYINPUT53), .A3(new_n1085), .A4(new_n1043), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1095));
  AOI211_X1 g670(.A(G171), .B(new_n1095), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1084), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1048), .A2(new_n725), .A3(new_n1051), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1966), .B1(new_n1045), .B2(new_n1043), .ZN(new_n1100));
  OAI21_X1  g675(.A(G8), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G286), .A2(G8), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT123), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1098), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1077), .A2(new_n756), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1048), .A2(new_n725), .A3(new_n1051), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1105), .A2(new_n1106), .B1(new_n1109), .B2(new_n1103), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1059), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT124), .B1(new_n1111), .B2(new_n1103), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1101), .A2(new_n1098), .A3(new_n1104), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(G2078), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1093), .B1(new_n1116), .B2(KEYINPUT53), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1088), .A2(G301), .A3(new_n1093), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT54), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1083), .A2(new_n1097), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n574), .B2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(new_n950), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1045), .A2(new_n1043), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1090), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1126), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1124), .A2(new_n1126), .A3(new_n1135), .A4(new_n1128), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1130), .A2(new_n1134), .A3(KEYINPUT122), .A4(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1090), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1058), .A2(new_n805), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1090), .A2(new_n1142), .B1(new_n805), .B2(new_n1058), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n608), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT60), .B(new_n883), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT58), .B(G1341), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1077), .A2(G1996), .B1(new_n1058), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n558), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT59), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1160), .B2(new_n1129), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1141), .A2(new_n1155), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n883), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1160), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1167), .A2(KEYINPUT120), .A3(new_n1129), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT120), .B1(new_n1167), .B2(new_n1129), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1121), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1052), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(new_n849), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1039), .B1(new_n1174), .B2(new_n1059), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1101), .A2(G286), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1057), .A3(new_n1075), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(G8), .B1(new_n1047), .B2(new_n1056), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1039), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1101), .A2(new_n1178), .A3(G286), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1057), .A3(new_n1075), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1112), .A2(KEYINPUT51), .A3(new_n1113), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1112), .B2(KEYINPUT51), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT62), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1076), .A2(new_n1082), .A3(new_n1118), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1110), .A2(new_n1190), .A3(new_n1114), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1057), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1071), .A2(new_n1072), .A3(new_n853), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1065), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1193), .A2(new_n1075), .B1(new_n1060), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1184), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1037), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1032), .A2(new_n1021), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT46), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n719), .A2(new_n1023), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1034), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1202), .B(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1024), .A2(new_n823), .A3(new_n820), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n803), .A2(new_n805), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1034), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1034), .A2(G1986), .A3(G290), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT48), .Z(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1033), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1205), .A2(new_n1206), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1198), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1216));
  INV_X1    g790(.A(G37), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n1216), .A2(new_n1005), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(KEYINPUT43), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1219), .A2(new_n1016), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n938), .A2(new_n944), .ZN(new_n1221));
  NOR2_X1   g795(.A1(G227), .A2(new_n461), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n657), .A2(new_n1222), .ZN(new_n1223));
  NOR3_X1   g797(.A1(new_n695), .A2(new_n696), .A3(new_n1223), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(G308));
  NAND3_X1  g799(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(G225));
endmodule


