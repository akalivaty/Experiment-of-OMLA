

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  NOR2_X1 U552 ( .A1(n533), .A2(n532), .ZN(n700) );
  XNOR2_X2 U553 ( .A(G2104), .B(KEYINPUT64), .ZN(n536) );
  BUF_X1 U554 ( .A(n737), .Z(n759) );
  AND2_X1 U555 ( .A1(n707), .A2(n706), .ZN(n713) );
  NAND2_X1 U556 ( .A1(n748), .A2(n747), .ZN(n758) );
  NAND2_X1 U557 ( .A1(n661), .A2(G56), .ZN(n599) );
  OR2_X1 U558 ( .A1(n713), .A2(n899), .ZN(n714) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n726) );
  NOR2_X1 U560 ( .A1(n775), .A2(n792), .ZN(n776) );
  INV_X1 U561 ( .A(KEYINPUT101), .ZN(n773) );
  AND2_X1 U562 ( .A1(n766), .A2(n765), .ZN(n767) );
  INV_X1 U563 ( .A(KEYINPUT104), .ZN(n795) );
  INV_X1 U564 ( .A(KEYINPUT23), .ZN(n521) );
  INV_X1 U565 ( .A(G2104), .ZN(n527) );
  INV_X1 U566 ( .A(KEYINPUT1), .ZN(n564) );
  NAND2_X1 U567 ( .A1(n610), .A2(n609), .ZN(n977) );
  BUF_X1 U568 ( .A(n700), .Z(G160) );
  AND2_X1 U569 ( .A1(n836), .A2(n826), .ZN(n517) );
  AND2_X1 U570 ( .A1(n830), .A2(n517), .ZN(n518) );
  AND2_X1 U571 ( .A1(n537), .A2(n536), .ZN(n519) );
  INV_X1 U572 ( .A(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U573 ( .A1(n751), .A2(n739), .ZN(n740) );
  XNOR2_X1 U574 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n730) );
  INV_X1 U575 ( .A(KEYINPUT100), .ZN(n749) );
  XNOR2_X1 U576 ( .A(n758), .B(n749), .ZN(n750) );
  INV_X1 U577 ( .A(KEYINPUT103), .ZN(n781) );
  INV_X1 U578 ( .A(KEYINPUT13), .ZN(n605) );
  NAND2_X1 U579 ( .A1(n527), .A2(n537), .ZN(n528) );
  INV_X1 U580 ( .A(KEYINPUT105), .ZN(n828) );
  XNOR2_X1 U581 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X1 U582 ( .A1(n608), .A2(n607), .ZN(n610) );
  BUF_X1 U583 ( .A(n701), .Z(G164) );
  INV_X1 U584 ( .A(G2105), .ZN(n537) );
  AND2_X1 U585 ( .A1(n537), .A2(G101), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n520), .A2(n536), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n553) );
  NAND2_X1 U589 ( .A1(n553), .A2(G125), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n526) );
  INV_X1 U591 ( .A(KEYINPUT65), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n533) );
  XNOR2_X2 U593 ( .A(n528), .B(KEYINPUT17), .ZN(n880) );
  NAND2_X1 U594 ( .A1(G137), .A2(n880), .ZN(n531) );
  NAND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U596 ( .A(KEYINPUT66), .B(n529), .Z(n884) );
  NAND2_X1 U597 ( .A1(G113), .A2(n884), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U599 ( .A1(G126), .A2(n553), .ZN(n535) );
  NAND2_X1 U600 ( .A1(G114), .A2(n884), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n541) );
  NAND2_X1 U602 ( .A1(G138), .A2(n880), .ZN(n539) );
  NAND2_X1 U603 ( .A1(G102), .A2(n519), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n701) );
  XNOR2_X1 U606 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U607 ( .A(G2451), .B(G2435), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n543) );
  XNOR2_X1 U609 ( .A(G2454), .B(G2430), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U611 ( .A(G2446), .B(G2438), .Z(n545) );
  XNOR2_X1 U612 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(n547), .B(n546), .Z(n549) );
  XNOR2_X1 U615 ( .A(G2443), .B(G2427), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U618 ( .A1(n552), .A2(G14), .ZN(G401) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U620 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n555) );
  BUF_X1 U621 ( .A(n553), .Z(n883) );
  NAND2_X1 U622 ( .A1(G123), .A2(n883), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G135), .A2(n880), .ZN(n557) );
  NAND2_X1 U625 ( .A1(G111), .A2(n884), .ZN(n556) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n519), .A2(G99), .ZN(n558) );
  XOR2_X1 U628 ( .A(KEYINPUT80), .B(n558), .Z(n559) );
  NOR2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n1008) );
  XNOR2_X1 U631 ( .A(G2096), .B(n1008), .ZN(n563) );
  OR2_X1 U632 ( .A1(G2100), .A2(n563), .ZN(G156) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  INV_X1 U635 ( .A(G69), .ZN(G235) );
  INV_X1 U636 ( .A(G108), .ZN(G238) );
  INV_X1 U637 ( .A(G120), .ZN(G236) );
  NOR2_X4 U638 ( .A1(G651), .A2(n639), .ZN(n669) );
  NAND2_X1 U639 ( .A1(G52), .A2(n669), .ZN(n567) );
  INV_X1 U640 ( .A(G651), .ZN(n569) );
  NOR2_X1 U641 ( .A1(G543), .A2(n569), .ZN(n565) );
  XNOR2_X2 U642 ( .A(n565), .B(n564), .ZN(n661) );
  NAND2_X1 U643 ( .A1(G64), .A2(n661), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U645 ( .A(KEYINPUT68), .B(n568), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n574) );
  NOR2_X2 U647 ( .A1(n639), .A2(n569), .ZN(n665) );
  NAND2_X1 U648 ( .A1(n665), .A2(G77), .ZN(n572) );
  NOR2_X1 U649 ( .A1(G651), .A2(G543), .ZN(n600) );
  BUF_X1 U650 ( .A(n600), .Z(n655) );
  NAND2_X1 U651 ( .A1(n655), .A2(G90), .ZN(n570) );
  XOR2_X1 U652 ( .A(KEYINPUT69), .B(n570), .Z(n571) );
  NAND2_X1 U653 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U654 ( .A(n574), .B(n573), .Z(n575) );
  NOR2_X1 U655 ( .A1(n576), .A2(n575), .ZN(G171) );
  NAND2_X1 U656 ( .A1(n655), .A2(G89), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n577), .B(KEYINPUT4), .ZN(n579) );
  NAND2_X1 U658 ( .A1(G76), .A2(n665), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n580), .B(KEYINPUT5), .ZN(n585) );
  NAND2_X1 U661 ( .A1(G51), .A2(n669), .ZN(n582) );
  NAND2_X1 U662 ( .A1(G63), .A2(n661), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U664 ( .A(KEYINPUT6), .B(n583), .Z(n584) );
  NAND2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U666 ( .A(n586), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U667 ( .A1(n661), .A2(G65), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G91), .A2(n655), .ZN(n588) );
  NAND2_X1 U669 ( .A1(G78), .A2(n665), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U671 ( .A1(G53), .A2(n669), .ZN(n589) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n589), .ZN(n590) );
  NOR2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U675 ( .A(n594), .B(KEYINPUT72), .ZN(G299) );
  XNOR2_X1 U676 ( .A(G168), .B(KEYINPUT8), .ZN(n595) );
  XNOR2_X1 U677 ( .A(n595), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U678 ( .A1(G7), .A2(G661), .ZN(n596) );
  XNOR2_X1 U679 ( .A(n596), .B(KEYINPUT10), .ZN(n597) );
  XNOR2_X1 U680 ( .A(KEYINPUT74), .B(n597), .ZN(G223) );
  INV_X1 U681 ( .A(G223), .ZN(n846) );
  NAND2_X1 U682 ( .A1(n846), .A2(G567), .ZN(n598) );
  XOR2_X1 U683 ( .A(KEYINPUT11), .B(n598), .Z(G234) );
  XOR2_X1 U684 ( .A(KEYINPUT14), .B(n599), .Z(n608) );
  NAND2_X1 U685 ( .A1(G81), .A2(n600), .ZN(n601) );
  XOR2_X1 U686 ( .A(KEYINPUT12), .B(n601), .Z(n602) );
  XNOR2_X1 U687 ( .A(n602), .B(KEYINPUT75), .ZN(n604) );
  NAND2_X1 U688 ( .A1(G68), .A2(n665), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n669), .A2(G43), .ZN(n609) );
  INV_X1 U691 ( .A(G860), .ZN(n624) );
  OR2_X1 U692 ( .A1(n977), .A2(n624), .ZN(G153) );
  INV_X1 U693 ( .A(G171), .ZN(G301) );
  NAND2_X1 U694 ( .A1(G868), .A2(G301), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G79), .A2(n665), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G66), .A2(n661), .ZN(n612) );
  NAND2_X1 U697 ( .A1(G92), .A2(n655), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n669), .A2(G54), .ZN(n613) );
  XOR2_X1 U700 ( .A(KEYINPUT76), .B(n613), .Z(n614) );
  NOR2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X2 U703 ( .A(n618), .B(KEYINPUT15), .ZN(n899) );
  INV_X1 U704 ( .A(n899), .ZN(n980) );
  INV_X1 U705 ( .A(G868), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n980), .A2(n621), .ZN(n619) );
  NAND2_X1 U707 ( .A1(n620), .A2(n619), .ZN(G284) );
  NOR2_X1 U708 ( .A1(G286), .A2(n621), .ZN(n623) );
  NOR2_X1 U709 ( .A1(G299), .A2(G868), .ZN(n622) );
  NOR2_X1 U710 ( .A1(n623), .A2(n622), .ZN(G297) );
  NAND2_X1 U711 ( .A1(n624), .A2(G559), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n625), .A2(n899), .ZN(n626) );
  XNOR2_X1 U713 ( .A(n626), .B(KEYINPUT16), .ZN(n627) );
  XNOR2_X1 U714 ( .A(KEYINPUT78), .B(n627), .ZN(G148) );
  NOR2_X1 U715 ( .A1(G868), .A2(n977), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n899), .A2(G868), .ZN(n628) );
  NOR2_X1 U717 ( .A1(G559), .A2(n628), .ZN(n629) );
  NOR2_X1 U718 ( .A1(n630), .A2(n629), .ZN(G282) );
  NAND2_X1 U719 ( .A1(G559), .A2(n899), .ZN(n631) );
  XNOR2_X1 U720 ( .A(n631), .B(n977), .ZN(n678) );
  NOR2_X1 U721 ( .A1(n678), .A2(G860), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G67), .A2(n661), .ZN(n633) );
  NAND2_X1 U723 ( .A1(G93), .A2(n655), .ZN(n632) );
  NAND2_X1 U724 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U725 ( .A1(G55), .A2(n669), .ZN(n635) );
  NAND2_X1 U726 ( .A1(G80), .A2(n665), .ZN(n634) );
  NAND2_X1 U727 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U728 ( .A1(n637), .A2(n636), .ZN(n681) );
  XNOR2_X1 U729 ( .A(n638), .B(n681), .ZN(G145) );
  NAND2_X1 U730 ( .A1(G49), .A2(n669), .ZN(n641) );
  NAND2_X1 U731 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U732 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U733 ( .A1(n661), .A2(n642), .ZN(n645) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n643) );
  XOR2_X1 U735 ( .A(KEYINPUT81), .B(n643), .Z(n644) );
  NAND2_X1 U736 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G47), .A2(n669), .ZN(n647) );
  NAND2_X1 U738 ( .A1(G60), .A2(n661), .ZN(n646) );
  NAND2_X1 U739 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U740 ( .A(KEYINPUT67), .B(n648), .ZN(n652) );
  NAND2_X1 U741 ( .A1(G85), .A2(n655), .ZN(n650) );
  NAND2_X1 U742 ( .A1(G72), .A2(n665), .ZN(n649) );
  AND2_X1 U743 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U744 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U745 ( .A1(G50), .A2(n669), .ZN(n654) );
  NAND2_X1 U746 ( .A1(G75), .A2(n665), .ZN(n653) );
  NAND2_X1 U747 ( .A1(n654), .A2(n653), .ZN(n659) );
  NAND2_X1 U748 ( .A1(G62), .A2(n661), .ZN(n657) );
  NAND2_X1 U749 ( .A1(G88), .A2(n655), .ZN(n656) );
  NAND2_X1 U750 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U751 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U752 ( .A(n660), .B(KEYINPUT83), .ZN(G303) );
  INV_X1 U753 ( .A(G303), .ZN(G166) );
  NAND2_X1 U754 ( .A1(G61), .A2(n661), .ZN(n663) );
  NAND2_X1 U755 ( .A1(G86), .A2(n655), .ZN(n662) );
  NAND2_X1 U756 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U757 ( .A(KEYINPUT82), .B(n664), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n665), .A2(G73), .ZN(n666) );
  XOR2_X1 U759 ( .A(KEYINPUT2), .B(n666), .Z(n667) );
  NOR2_X1 U760 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n669), .A2(G48), .ZN(n670) );
  NAND2_X1 U762 ( .A1(n671), .A2(n670), .ZN(G305) );
  XNOR2_X1 U763 ( .A(KEYINPUT84), .B(G288), .ZN(n672) );
  XNOR2_X1 U764 ( .A(n672), .B(G290), .ZN(n673) );
  XOR2_X1 U765 ( .A(n673), .B(KEYINPUT19), .Z(n675) );
  XNOR2_X1 U766 ( .A(G166), .B(n681), .ZN(n674) );
  XNOR2_X1 U767 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U768 ( .A(n676), .B(G305), .Z(n677) );
  XNOR2_X1 U769 ( .A(G299), .B(n677), .ZN(n895) );
  XNOR2_X1 U770 ( .A(KEYINPUT85), .B(n678), .ZN(n679) );
  XNOR2_X1 U771 ( .A(n895), .B(n679), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n680), .A2(G868), .ZN(n683) );
  OR2_X1 U773 ( .A1(G868), .A2(n681), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n683), .A2(n682), .ZN(G295) );
  NAND2_X1 U775 ( .A1(G2084), .A2(G2078), .ZN(n684) );
  XOR2_X1 U776 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U777 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U778 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U779 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U780 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U781 ( .A1(G237), .A2(G236), .ZN(n689) );
  NOR2_X1 U782 ( .A1(G238), .A2(G235), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U784 ( .A(KEYINPUT86), .B(n690), .ZN(n852) );
  NAND2_X1 U785 ( .A1(n852), .A2(G567), .ZN(n691) );
  XNOR2_X1 U786 ( .A(n691), .B(KEYINPUT87), .ZN(n696) );
  NOR2_X1 U787 ( .A1(G220), .A2(G219), .ZN(n692) );
  XNOR2_X1 U788 ( .A(KEYINPUT22), .B(n692), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n693), .A2(G96), .ZN(n694) );
  OR2_X1 U790 ( .A1(G218), .A2(n694), .ZN(n851) );
  AND2_X1 U791 ( .A1(G2106), .A2(n851), .ZN(n695) );
  NOR2_X1 U792 ( .A1(n696), .A2(n695), .ZN(G319) );
  NAND2_X1 U793 ( .A1(G483), .A2(G661), .ZN(n698) );
  INV_X1 U794 ( .A(G319), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U796 ( .A(n699), .B(KEYINPUT88), .ZN(n849) );
  NAND2_X1 U797 ( .A1(G36), .A2(n849), .ZN(G176) );
  NAND2_X1 U798 ( .A1(n700), .A2(G40), .ZN(n815) );
  INV_X1 U799 ( .A(n815), .ZN(n702) );
  NOR2_X2 U800 ( .A1(n701), .A2(G1384), .ZN(n816) );
  NAND2_X2 U801 ( .A1(n702), .A2(n816), .ZN(n737) );
  NAND2_X1 U802 ( .A1(G8), .A2(n759), .ZN(n792) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n792), .ZN(n751) );
  INV_X1 U804 ( .A(G1996), .ZN(n929) );
  NOR2_X1 U805 ( .A1(n737), .A2(n929), .ZN(n704) );
  XNOR2_X1 U806 ( .A(n704), .B(n703), .ZN(n707) );
  AND2_X1 U807 ( .A1(n737), .A2(G1341), .ZN(n705) );
  NOR2_X1 U808 ( .A1(n705), .A2(n977), .ZN(n706) );
  NAND2_X1 U809 ( .A1(n713), .A2(n899), .ZN(n712) );
  AND2_X1 U810 ( .A1(n759), .A2(G1348), .ZN(n708) );
  XNOR2_X1 U811 ( .A(n708), .B(KEYINPUT97), .ZN(n710) );
  INV_X1 U812 ( .A(n737), .ZN(n732) );
  NAND2_X1 U813 ( .A1(n732), .A2(G2067), .ZN(n709) );
  NAND2_X1 U814 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U815 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U817 ( .A(n716), .B(KEYINPUT98), .ZN(n723) );
  INV_X1 U818 ( .A(G299), .ZN(n724) );
  INV_X1 U819 ( .A(n737), .ZN(n717) );
  NAND2_X1 U820 ( .A1(n717), .A2(G2072), .ZN(n718) );
  XNOR2_X1 U821 ( .A(n718), .B(KEYINPUT27), .ZN(n720) );
  XNOR2_X1 U822 ( .A(KEYINPUT95), .B(G1956), .ZN(n963) );
  NOR2_X1 U823 ( .A1(n963), .A2(n732), .ZN(n719) );
  NOR2_X1 U824 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U825 ( .A(KEYINPUT96), .B(n721), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n724), .A2(n725), .ZN(n722) );
  NAND2_X1 U827 ( .A1(n723), .A2(n722), .ZN(n729) );
  NOR2_X1 U828 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U829 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U831 ( .A(n731), .B(n730), .ZN(n736) );
  XOR2_X1 U832 ( .A(KEYINPUT25), .B(G2078), .Z(n934) );
  NOR2_X1 U833 ( .A1(n934), .A2(n759), .ZN(n734) );
  NOR2_X1 U834 ( .A1(n732), .A2(G1961), .ZN(n733) );
  NOR2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n743) );
  OR2_X1 U836 ( .A1(G301), .A2(n743), .ZN(n735) );
  NAND2_X1 U837 ( .A1(n736), .A2(n735), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n737), .A2(G2084), .ZN(n738) );
  XNOR2_X1 U839 ( .A(n738), .B(KEYINPUT93), .ZN(n752) );
  NAND2_X1 U840 ( .A1(G8), .A2(n752), .ZN(n739) );
  XNOR2_X1 U841 ( .A(n740), .B(KEYINPUT30), .ZN(n742) );
  INV_X1 U842 ( .A(G168), .ZN(n741) );
  NAND2_X1 U843 ( .A1(n742), .A2(n741), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n743), .A2(G301), .ZN(n744) );
  NAND2_X1 U845 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U846 ( .A(n746), .B(KEYINPUT31), .ZN(n747) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n756) );
  INV_X1 U848 ( .A(n752), .ZN(n753) );
  NAND2_X1 U849 ( .A1(n753), .A2(G8), .ZN(n754) );
  XNOR2_X1 U850 ( .A(n754), .B(KEYINPUT94), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n756), .A2(n755), .ZN(n769) );
  AND2_X1 U852 ( .A1(G286), .A2(G8), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n766) );
  INV_X1 U854 ( .A(G8), .ZN(n764) );
  NOR2_X1 U855 ( .A1(G1971), .A2(n792), .ZN(n761) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U857 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n762), .A2(G303), .ZN(n763) );
  OR2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U860 ( .A(n767), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n786) );
  NOR2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U864 ( .A1(n983), .A2(n770), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n786), .A2(n771), .ZN(n772) );
  NAND2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NAND2_X1 U867 ( .A1(n772), .A2(n986), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(n773), .ZN(n775) );
  NOR2_X1 U869 ( .A1(n776), .A2(KEYINPUT33), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n983), .A2(KEYINPUT33), .ZN(n777) );
  XNOR2_X1 U871 ( .A(KEYINPUT102), .B(n777), .ZN(n778) );
  NOR2_X1 U872 ( .A1(n778), .A2(n792), .ZN(n779) );
  NOR2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n782) );
  XNOR2_X1 U874 ( .A(n782), .B(n781), .ZN(n783) );
  XOR2_X1 U875 ( .A(G1981), .B(G305), .Z(n995) );
  NAND2_X1 U876 ( .A1(n783), .A2(n995), .ZN(n789) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U878 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n787), .A2(n792), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n794) );
  NOR2_X1 U882 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U883 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  NOR2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(n795), .ZN(n827) );
  NAND2_X1 U887 ( .A1(G141), .A2(n880), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G117), .A2(n884), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n519), .A2(G105), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n883), .A2(G129), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n875) );
  NAND2_X1 U895 ( .A1(n875), .A2(G1996), .ZN(n813) );
  XNOR2_X1 U896 ( .A(KEYINPUT90), .B(G1991), .ZN(n933) );
  NAND2_X1 U897 ( .A1(G131), .A2(n880), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G107), .A2(n884), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G95), .A2(n519), .ZN(n806) );
  XNOR2_X1 U901 ( .A(KEYINPUT89), .B(n806), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n883), .A2(G119), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n890) );
  NAND2_X1 U905 ( .A1(n933), .A2(n890), .ZN(n811) );
  XOR2_X1 U906 ( .A(KEYINPUT91), .B(n811), .Z(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT92), .ZN(n1024) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n841) );
  NAND2_X1 U910 ( .A1(n1024), .A2(n841), .ZN(n830) );
  NAND2_X1 U911 ( .A1(G104), .A2(n519), .ZN(n818) );
  NAND2_X1 U912 ( .A1(G140), .A2(n880), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U914 ( .A(KEYINPUT34), .B(n819), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G128), .A2(n883), .ZN(n821) );
  NAND2_X1 U916 ( .A1(G116), .A2(n884), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U918 ( .A(KEYINPUT35), .B(n822), .Z(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT36), .B(n825), .ZN(n877) );
  XNOR2_X1 U921 ( .A(G2067), .B(KEYINPUT37), .ZN(n838) );
  NOR2_X1 U922 ( .A1(n877), .A2(n838), .ZN(n1007) );
  NAND2_X1 U923 ( .A1(n841), .A2(n1007), .ZN(n836) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U925 ( .A1(n841), .A2(n982), .ZN(n826) );
  NAND2_X1 U926 ( .A1(n827), .A2(n518), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n844) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n875), .ZN(n1003) );
  INV_X1 U929 ( .A(n830), .ZN(n833) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n831) );
  NOR2_X1 U931 ( .A1(n933), .A2(n890), .ZN(n1011) );
  NOR2_X1 U932 ( .A1(n831), .A2(n1011), .ZN(n832) );
  NOR2_X1 U933 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U934 ( .A1(n1003), .A2(n834), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U937 ( .A1(n877), .A2(n838), .ZN(n1012) );
  NAND2_X1 U938 ( .A1(n839), .A2(n1012), .ZN(n840) );
  NAND2_X1 U939 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U940 ( .A(KEYINPUT106), .B(n842), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U945 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(KEYINPUT109), .B(n850), .Z(G188) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  NOR2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT110), .B(n853), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  NAND2_X1 U954 ( .A1(G100), .A2(n519), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G112), .A2(n884), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n883), .A2(G124), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G136), .A2(n880), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U963 ( .A(G164), .B(KEYINPUT112), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT113), .B(n863), .ZN(n874) );
  NAND2_X1 U966 ( .A1(G130), .A2(n883), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G118), .A2(n884), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G106), .A2(n519), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G142), .A2(n880), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(KEYINPUT45), .B(n868), .ZN(n869) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n869), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n1008), .B(n872), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U979 ( .A(G162), .B(n879), .ZN(n892) );
  NAND2_X1 U980 ( .A1(G103), .A2(n519), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G127), .A2(n883), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G115), .A2(n884), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n1014) );
  XNOR2_X1 U988 ( .A(n890), .B(n1014), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(G160), .B(n893), .Z(n894) );
  NOR2_X1 U991 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U992 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n977), .B(n895), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n898), .B(G286), .Z(n901) );
  XNOR2_X1 U996 ( .A(n899), .B(G171), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2100), .B(G2096), .Z(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT42), .B(G2678), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1002 ( .A(KEYINPUT43), .B(G2090), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G2072), .B(G2067), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G2084), .B(G2078), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(G227) );
  XOR2_X1 U1008 ( .A(G1981), .B(G1961), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G1956), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1011 ( .A(n913), .B(KEYINPUT41), .Z(n915) );
  XNOR2_X1 U1012 ( .A(G1996), .B(G1991), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n919) );
  XOR2_X1 U1014 ( .A(G2474), .B(G1986), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G1971), .B(G1976), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(G229) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT117), .B(n920), .Z(n926) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n921), .Z(n922) );
  NAND2_X1 U1022 ( .A1(G319), .A2(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(G401), .A2(n923), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1027 ( .A(KEYINPUT121), .B(G34), .Z(n928) );
  XNOR2_X1 U1028 ( .A(G2084), .B(KEYINPUT54), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(n928), .B(n927), .ZN(n946) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G35), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(G32), .B(n929), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n930), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G2072), .B(G33), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n933), .B(G25), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G27), .B(n934), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1043 ( .A(KEYINPUT120), .B(n944), .Z(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(KEYINPUT55), .B(n947), .ZN(n949) );
  INV_X1 U1046 ( .A(G29), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n950), .A2(G11), .ZN(n951) );
  XOR2_X1 U1049 ( .A(KEYINPUT122), .B(n951), .Z(n1034) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G22), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G24), .B(G1986), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1053 ( .A(G1976), .B(G23), .Z(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n957) );
  XOR2_X1 U1055 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n956) );
  XNOR2_X1 U1056 ( .A(n957), .B(n956), .ZN(n971) );
  XNOR2_X1 U1057 ( .A(G1348), .B(KEYINPUT59), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(n958), .B(G4), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G1341), .B(G19), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(G6), .B(G1981), .ZN(n959) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n963), .ZN(n964) );
  XNOR2_X1 U1064 ( .A(G20), .B(n964), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1066 ( .A(KEYINPUT60), .B(n967), .Z(n969) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G21), .ZN(n968) );
  NOR2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G5), .B(G1961), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1072 ( .A(KEYINPUT61), .B(n974), .Z(n975) );
  NOR2_X1 U1073 ( .A1(G16), .A2(n975), .ZN(n976) );
  XOR2_X1 U1074 ( .A(KEYINPUT127), .B(n976), .Z(n1032) );
  XNOR2_X1 U1075 ( .A(KEYINPUT56), .B(G16), .ZN(n1001) );
  XOR2_X1 U1076 ( .A(n977), .B(G1341), .Z(n979) );
  XNOR2_X1 U1077 ( .A(G171), .B(G1961), .ZN(n978) );
  NAND2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n980), .ZN(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n991) );
  XOR2_X1 U1081 ( .A(n983), .B(KEYINPUT123), .Z(n985) );
  XOR2_X1 U1082 ( .A(G166), .B(G1971), .Z(n984) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n988) );
  NOR2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT124), .B(n994), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(KEYINPUT57), .B(n997), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1030) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1004), .Z(n1005) );
  XOR2_X1 U1098 ( .A(KEYINPUT118), .B(n1005), .Z(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1022) );
  XNOR2_X1 U1100 ( .A(G160), .B(G2084), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(G2072), .B(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(G164), .B(G2078), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1107 ( .A(KEYINPUT50), .B(n1017), .Z(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT119), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1025), .ZN(n1027) );
  INV_X1 U1113 ( .A(KEYINPUT55), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(G29), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

