//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT66), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n462), .A2(new_n463), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n462), .B2(new_n463), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n463), .C2(new_n462), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g077(.A(G651), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT68), .A2(G88), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT68), .A2(G88), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n503), .A2(new_n505), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n511), .B2(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n503), .A2(new_n513), .A3(G50), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n510), .B(new_n514), .C1(new_n515), .C2(new_n504), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  XNOR2_X1  g092(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n512), .B1(new_n518), .B2(G651), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT69), .B(G51), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n511), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n504), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n505), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n523), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT70), .B1(new_n521), .B2(new_n522), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n504), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n519), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n533), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n533), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n530), .A2(new_n531), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n503), .A2(new_n513), .A3(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT72), .B1(new_n560), .B2(new_n504), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n547), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT71), .B1(new_n529), .B2(new_n532), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n503), .A2(new_n569), .A3(new_n505), .A4(new_n509), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G91), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n559), .A2(new_n567), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  OR2_X1    g148(.A1(new_n509), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n519), .B2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n568), .A2(G87), .A3(new_n570), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n578));
  OAI21_X1  g153(.A(G61), .B1(new_n530), .B2(new_n531), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(G651), .ZN(new_n582));
  AOI211_X1 g157(.A(KEYINPUT73), .B(new_n504), .C1(new_n579), .C2(new_n580), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n519), .A2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n568), .A2(G86), .A3(new_n570), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n584), .A2(new_n589), .A3(new_n585), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n533), .A2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n519), .A2(G47), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n504), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n519), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n504), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n568), .A2(new_n570), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  XNOR2_X1  g185(.A(G280), .B(KEYINPUT75), .ZN(G297));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n551), .A2(new_n608), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n612), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g193(.A(KEYINPUT3), .B(G2104), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n465), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G123), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(G156));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n636), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(new_n648), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT76), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n650), .A3(new_n648), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n650), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n659), .B1(new_n649), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  AOI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT77), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(G229));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n684));
  NAND2_X1  g259(.A1(G103), .A2(G2104), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G2105), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n479), .A2(G139), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n619), .A2(G127), .ZN(new_n689));
  NAND2_X1  g264(.A1(G115), .A2(G2104), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n461), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n688), .B1(KEYINPUT82), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(KEYINPUT82), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G33), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2072), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(G34), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT78), .B(G29), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(G34), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n476), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G2084), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n699), .A2(G35), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G162), .B2(new_n699), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT87), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G2090), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n705), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n696), .B(new_n713), .C1(new_n712), .C2(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n552), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G16), .B2(G19), .ZN(new_n716));
  INV_X1    g291(.A(G1341), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n479), .A2(G140), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n481), .A2(G128), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n461), .A2(G116), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n700), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G5), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G301), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(new_n717), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n718), .A2(new_n729), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT31), .B(G11), .Z(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT85), .B(G28), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n630), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n703), .A2(G32), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n481), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n742), .B1(new_n743), .B2(new_n700), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n699), .A2(G27), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n699), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n732), .A2(new_n733), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n753), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  NOR2_X1   g335(.A1(G4), .A2(G16), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n605), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n736), .B(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n730), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n730), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT84), .B(G1966), .Z(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G1348), .B2(new_n762), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n730), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT89), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n714), .A2(new_n764), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n730), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n730), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1971), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G23), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT80), .Z(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G288), .B2(new_n730), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(G6), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G305), .B2(new_n730), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT34), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n793), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n700), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n479), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n481), .A2(G119), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n461), .A2(G107), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n799), .B1(new_n808), .B2(new_n699), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1986), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n796), .A2(new_n798), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT81), .B(KEYINPUT36), .Z(new_n817));
  AOI21_X1  g392(.A(new_n778), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n819));
  INV_X1    g394(.A(new_n816), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n820), .A2(KEYINPUT81), .A3(KEYINPUT36), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n819), .B1(new_n818), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n818), .A2(new_n821), .ZN(G150));
  NAND2_X1  g400(.A1(new_n533), .A2(G93), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT91), .B(G55), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n519), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT92), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n547), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n830), .A2(new_n832), .B1(G651), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT96), .B(G860), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n603), .A2(new_n604), .ZN(new_n841));
  INV_X1    g416(.A(new_n599), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n612), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n830), .A2(new_n832), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n835), .A2(G651), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n544), .A2(new_n550), .A3(new_n545), .A4(KEYINPUT93), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n551), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n551), .B2(new_n851), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n836), .A2(new_n857), .A3(new_n849), .A4(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n846), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n845), .A2(new_n858), .A3(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT95), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n860), .A2(new_n864), .A3(new_n865), .A4(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n838), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n840), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT97), .ZN(G145));
  NAND2_X1  g445(.A1(new_n497), .A2(new_n499), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n490), .A2(new_n492), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n723), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n749), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(new_n694), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT100), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n694), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n806), .A2(KEYINPUT102), .A3(new_n807), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n806), .B2(new_n807), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n621), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n479), .A2(G142), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n481), .A2(G130), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n808), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n621), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n884), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n887), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n887), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n883), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT103), .A3(new_n898), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n879), .A2(new_n882), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n476), .B(KEYINPUT98), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G162), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n743), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n879), .A2(new_n882), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n899), .A2(new_n900), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n904), .B(new_n908), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n901), .A2(new_n903), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n904), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n907), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n914), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT40), .B1(new_n914), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G395));
  OAI21_X1  g496(.A(KEYINPUT108), .B1(new_n836), .B2(G868), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n859), .A2(new_n616), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n856), .A2(new_n615), .A3(new_n858), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n843), .A2(G299), .ZN(new_n926));
  INV_X1    g501(.A(G299), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n605), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT41), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n925), .A2(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT107), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(G288), .B(G290), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n588), .A2(G303), .A3(new_n590), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G303), .B1(new_n588), .B2(new_n590), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n943), .A3(new_n945), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT106), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT106), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n950), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n608), .B1(new_n942), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n939), .A2(new_n941), .A3(new_n955), .A4(new_n958), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n922), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  INV_X1    g538(.A(new_n941), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n935), .A2(new_n940), .A3(KEYINPUT107), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n959), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n963), .A2(new_n966), .A3(G868), .A4(new_n961), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n962), .A2(new_n967), .ZN(G295));
  NOR2_X1   g543(.A1(new_n962), .A2(new_n967), .ZN(G331));
  XOR2_X1   g544(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n856), .A2(G301), .A3(new_n858), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G301), .B1(new_n856), .B2(new_n858), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(G286), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n859), .A2(G171), .ZN(new_n976));
  AOI21_X1  g551(.A(G168), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n934), .B(new_n933), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G286), .B1(new_n973), .B2(new_n974), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(G168), .A3(new_n972), .ZN(new_n980));
  INV_X1    g555(.A(new_n929), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n953), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G37), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n953), .B1(new_n978), .B2(new_n982), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n971), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n979), .A2(new_n980), .A3(new_n988), .A4(new_n981), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n979), .A2(new_n980), .B1(new_n932), .B2(new_n930), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n954), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n984), .A3(new_n983), .A4(new_n970), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n984), .A3(new_n983), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  INV_X1    g573(.A(new_n986), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(new_n984), .A3(new_n983), .A4(new_n970), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  INV_X1    g578(.A(new_n499), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n498), .B1(new_n619), .B2(new_n495), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n874), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n619), .A2(new_n491), .B1(new_n1008), .B2(new_n489), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n873), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT112), .B(G40), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n474), .B2(G2105), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n469), .A3(new_n470), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n723), .B(G2067), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT114), .Z(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(G1996), .A3(new_n749), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1017), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(G1996), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n749), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n806), .A2(new_n810), .A3(new_n807), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n810), .B1(new_n806), .B2(new_n807), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1017), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G290), .B(G1986), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1017), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT127), .ZN(new_n1033));
  AND3_X1   g608(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT45), .B(new_n1003), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1015), .A2(new_n470), .A3(new_n469), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT115), .B(G1971), .Z(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1384), .B1(new_n871), .B2(new_n1009), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1016), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT116), .B(G8), .Z(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1037), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n875), .A2(new_n1044), .A3(new_n1003), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1048), .A3(new_n1039), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1043), .B2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1053), .A2(KEYINPUT119), .B1(new_n1037), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1051), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n1037), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT73), .B1(new_n1064), .B2(new_n504), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n581), .A2(new_n578), .A3(G651), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1981), .B1(new_n519), .B2(G48), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n586), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n584), .A2(new_n1070), .A3(new_n586), .A4(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n533), .A2(G86), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n585), .C1(new_n504), .C2(new_n1064), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G1981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1072), .A2(new_n1078), .A3(KEYINPUT49), .A4(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT49), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1011), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1039), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1052), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n575), .A2(new_n576), .A3(G1976), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1052), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(new_n1052), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1033), .B1(new_n1063), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1009), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1044), .A3(new_n1003), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1039), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1044), .B1(new_n875), .B2(new_n1003), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1101), .A2(new_n1048), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT119), .B(new_n1036), .C1(new_n1102), .C2(new_n1051), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1058), .A2(new_n1037), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1062), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1093), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT127), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1055), .A2(new_n1039), .A3(new_n1056), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(G2084), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1016), .B1(KEYINPUT45), .B2(new_n1045), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n768), .B1(new_n1110), .B2(new_n1013), .ZN(new_n1111));
  OAI21_X1  g686(.A(G8), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G286), .A2(new_n1052), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1052), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1114), .B(KEYINPUT51), .C1(G168), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(new_n1113), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1108), .A2(KEYINPUT124), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1055), .A2(new_n1121), .A3(new_n1039), .A4(new_n1056), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n733), .A3(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1110), .A2(new_n1013), .A3(KEYINPUT53), .A4(new_n756), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1041), .B2(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1096), .A2(new_n1107), .B1(new_n1119), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(G301), .B(KEYINPUT54), .Z(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n756), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1132));
  NAND4_X1  g707(.A1(G160), .A2(new_n1013), .A3(new_n1038), .A4(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1123), .A2(new_n1126), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1134), .B2(new_n1130), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n927), .B2(KEYINPUT122), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  NAND3_X1  g713(.A1(G299), .A2(new_n1138), .A3(KEYINPUT57), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1956), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(G2072), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1038), .A2(new_n1040), .A3(new_n1039), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1140), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1137), .A2(new_n1146), .A3(new_n1142), .A4(new_n1139), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT126), .B(G1996), .Z(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1041), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n552), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n552), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1150), .A2(new_n1151), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1120), .A2(new_n760), .A3(new_n1122), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1082), .A2(new_n728), .A3(new_n1039), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(KEYINPUT60), .A3(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n605), .A3(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(new_n605), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1147), .A2(KEYINPUT125), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1142), .A2(new_n1170), .A3(new_n1146), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1171), .A3(new_n1140), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1160), .A2(new_n1167), .A3(new_n1168), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1163), .A2(new_n605), .A3(new_n1149), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1175), .A2(new_n1172), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1135), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1127), .A2(G171), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1119), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(KEYINPUT62), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1129), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1086), .A2(new_n1182), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1183), .A2(new_n1084), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1115), .A2(G286), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1106), .A2(new_n1059), .A3(new_n1062), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1105), .A2(new_n1189), .A3(new_n1106), .A4(new_n1185), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1058), .A2(new_n1037), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1192), .A2(G286), .A3(new_n1115), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1193), .A2(new_n1106), .A3(KEYINPUT63), .A4(new_n1104), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1184), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1181), .B1(new_n1195), .B2(KEYINPUT121), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1197), .B(new_n1184), .C1(new_n1191), .C2(new_n1194), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1032), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1024), .A2(KEYINPUT46), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1024), .A2(KEYINPUT46), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1018), .A2(new_n749), .ZN(new_n1202));
  AOI22_X1  g777(.A1(new_n1200), .A2(new_n1201), .B1(new_n1017), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n723), .A2(G2067), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1023), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1023), .A2(G1986), .A3(G290), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT48), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1030), .A2(new_n1209), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1204), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1199), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g787(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n681), .A2(new_n682), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1215), .B1(new_n914), .B2(new_n918), .ZN(new_n1216));
  AND2_X1   g790(.A1(new_n1216), .A2(new_n994), .ZN(G308));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n994), .ZN(G225));
endmodule


