//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000;
  XNOR2_X1  g000(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT90), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G141gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G169gat), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT12), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G15gat), .B(G22gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G1gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT91), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(G8gat), .B1(new_n216), .B2(KEYINPUT92), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n214), .B(new_n211), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI221_X1 g020(.A(new_n216), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n218), .C2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G29gat), .A2(G36gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230));
  NAND2_X1  g029(.A1(G43gat), .A2(G50gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G29gat), .A2(G36gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n231), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT15), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n232), .A2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(KEYINPUT15), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(new_n226), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n223), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT13), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n221), .A2(new_n222), .A3(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n238), .A2(new_n226), .A3(new_n232), .A4(new_n233), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n238), .B1(new_n237), .B2(new_n226), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT17), .A3(new_n239), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT93), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n223), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n221), .A2(KEYINPUT93), .A3(new_n222), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n248), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT94), .B1(new_n258), .B2(new_n242), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n246), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n223), .A2(new_n255), .ZN(new_n262));
  INV_X1    g061(.A(new_n254), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(new_n242), .A3(new_n247), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT18), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n209), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n245), .B1(new_n267), .B2(KEYINPUT18), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n260), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n208), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G113gat), .B2(G120gat), .ZN(new_n277));
  AND2_X1   g076(.A1(G113gat), .A2(G120gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  INV_X1    g079(.A(G127gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n275), .B(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(G134gat), .A3(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT27), .B(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT28), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT27), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n294));
  AOI21_X1  g093(.A(G190gat), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n295), .B2(KEYINPUT28), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT66), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n298), .A2(new_n303), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n299), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n291), .A2(new_n292), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n307), .B1(new_n319), .B2(new_n289), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n308), .B(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n318), .B1(new_n323), .B2(new_n317), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n287), .B1(new_n305), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G227gat), .ZN(new_n326));
  INV_X1    g125(.A(G233gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n280), .A2(G134gat), .A3(new_n282), .ZN(new_n329));
  AOI21_X1  g128(.A(G134gat), .B1(new_n280), .B2(new_n282), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n310), .A2(new_n315), .A3(KEYINPUT25), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n308), .B(KEYINPUT64), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT65), .B(G183gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n306), .B1(new_n334), .B2(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n316), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n336), .B2(KEYINPUT25), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n296), .A2(new_n304), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n325), .A2(new_n328), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT68), .B(G71gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G99gat), .ZN(new_n345));
  XOR2_X1   g144(.A(G15gat), .B(G43gat), .Z(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n340), .B(KEYINPUT32), .C1(new_n342), .C2(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n339), .ZN(new_n352));
  INV_X1    g151(.A(new_n328), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n352), .A2(KEYINPUT34), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT34), .B1(new_n352), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT71), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n350), .A3(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n358), .A2(KEYINPUT71), .A3(new_n349), .A4(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n352), .A2(KEYINPUT34), .A3(new_n353), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT69), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n354), .B2(new_n355), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n351), .A2(new_n365), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n359), .A3(new_n371), .ZN(new_n372));
  MUX2_X1   g171(.A(new_n362), .B(new_n372), .S(KEYINPUT36), .Z(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G211gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT72), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G211gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT22), .B1(new_n381), .B2(G218gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n376), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT22), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT72), .B(G211gat), .ZN(new_n387));
  INV_X1    g186(.A(G218gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(new_n375), .A3(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT73), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n393));
  XNOR2_X1  g192(.A(G155gat), .B(G162gat), .ZN(new_n394));
  AND2_X1   g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  INV_X1    g201(.A(G141gat), .ZN(new_n403));
  INV_X1    g202(.A(G148gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n409), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT80), .B1(new_n409), .B2(KEYINPUT2), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n394), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n408), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n415), .B2(new_n398), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n409), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n407), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT81), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n393), .B(new_n400), .C1(new_n414), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n374), .B1(new_n392), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n400), .B1(new_n414), .B2(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT82), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n413), .B1(new_n408), .B2(new_n412), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n421), .A2(KEYINPUT81), .A3(new_n422), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n399), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT3), .B1(new_n391), .B2(new_n425), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n389), .A2(new_n438), .A3(new_n375), .A4(new_n383), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(new_n425), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n385), .A2(KEYINPUT85), .A3(new_n390), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n432), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n391), .B1(new_n424), .B2(new_n425), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT86), .B(new_n374), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n432), .B2(new_n393), .ZN(new_n447));
  OAI22_X1  g246(.A1(new_n447), .A2(new_n391), .B1(new_n442), .B2(new_n432), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT86), .B1(new_n448), .B2(new_n374), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n437), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G22gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n374), .B1(new_n443), .B2(new_n444), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n445), .ZN(new_n455));
  INV_X1    g254(.A(G22gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n437), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT31), .B(G50gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n451), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n451), .B2(new_n457), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n428), .B2(new_n331), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n287), .A3(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT3), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n287), .B1(new_n432), .B2(new_n393), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  OR3_X1    g270(.A1(new_n470), .A2(KEYINPUT39), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n432), .A2(new_n287), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n430), .A2(new_n431), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n433), .B1(new_n475), .B2(new_n400), .ZN(new_n476));
  AOI211_X1 g275(.A(KEYINPUT82), .B(new_n399), .C1(new_n430), .C2(new_n431), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(new_n331), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(KEYINPUT39), .C1(new_n471), .C2(new_n470), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n482));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G57gat), .B(G85gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND4_X1  g285(.A1(new_n472), .A2(new_n481), .A3(KEYINPUT40), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n471), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT5), .B1(new_n479), .B2(new_n471), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n488), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n466), .A3(new_n465), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n468), .B2(new_n469), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n490), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n486), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n472), .A2(new_n481), .A3(new_n486), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT74), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n305), .B2(new_n324), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT74), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n502), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT29), .B1(new_n337), .B2(new_n338), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n506), .A2(KEYINPUT75), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n392), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT29), .B1(new_n504), .B2(new_n505), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(new_n507), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT74), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT74), .B1(new_n337), .B2(new_n338), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n425), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT76), .A3(new_n502), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n507), .B1(new_n305), .B2(new_n324), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT77), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n514), .A2(new_n518), .A3(new_n391), .A4(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G36gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT78), .B(G8gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n511), .A2(new_n521), .A3(KEYINPUT30), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n521), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n525), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n463), .B1(new_n501), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n473), .B1(new_n435), .B2(new_n287), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(new_n488), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n468), .A2(new_n469), .ZN(new_n540));
  INV_X1    g339(.A(new_n467), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n492), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n486), .B1(new_n543), .B2(new_n490), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT6), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n539), .A2(new_n542), .B1(new_n470), .B2(new_n489), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT6), .B1(new_n547), .B2(new_n486), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n536), .A2(new_n546), .B1(new_n497), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n509), .A2(new_n510), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n514), .A2(new_n518), .A3(new_n520), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n550), .A2(new_n392), .B1(new_n551), .B2(new_n391), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT38), .B1(new_n552), .B2(KEYINPUT37), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n511), .A2(new_n521), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n525), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n511), .B2(new_n521), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT38), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n549), .A2(new_n558), .A3(new_n527), .A4(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n373), .B1(new_n534), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n536), .A2(new_n546), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n497), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n533), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n460), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n450), .A2(G22gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n456), .B1(new_n455), .B2(new_n437), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n451), .A2(new_n457), .A3(new_n460), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n569), .A2(KEYINPUT87), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT87), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n562), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n463), .B2(new_n372), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n369), .A2(new_n359), .A3(new_n371), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n570), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT88), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(KEYINPUT35), .A3(new_n565), .A4(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n545), .B1(new_n544), .B2(KEYINPUT6), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT6), .ZN(new_n583));
  NOR4_X1   g382(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n583), .A4(new_n486), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n564), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n533), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n362), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n274), .B1(new_n574), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI221_X1 g399(.A(new_n593), .B1(new_n598), .B2(new_n597), .C1(new_n594), .C2(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT20), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n607), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n602), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n223), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G183gat), .ZN(new_n616));
  INV_X1    g415(.A(G183gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n617), .A3(new_n223), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n607), .B(new_n609), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G211gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n623), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT8), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(KEYINPUT100), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(KEYINPUT100), .B2(new_n629), .ZN(new_n631));
  OR2_X1    g430(.A1(KEYINPUT101), .A2(G85gat), .ZN(new_n632));
  INV_X1    g431(.A(G92gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT101), .A2(G85gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G85gat), .A2(G92gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT7), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G99gat), .B(G106gat), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT102), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n642), .A3(new_n639), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n263), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G190gat), .B(G218gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n646), .A2(new_n240), .B1(KEYINPUT41), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n650), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n650), .A2(new_n654), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n651), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n656), .A3(new_n655), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n655), .A4(new_n661), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n655), .A3(new_n661), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n627), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(G230gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n327), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n602), .A2(new_n612), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n600), .B2(new_n601), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT10), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n645), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n641), .A2(new_n603), .A3(new_n644), .A4(new_n643), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n638), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n639), .ZN(new_n683));
  INV_X1    g482(.A(new_n639), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n638), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n602), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT10), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n675), .B1(new_n679), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n680), .A2(new_n674), .A3(new_n686), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G176gat), .ZN(new_n692));
  INV_X1    g491(.A(G204gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n690), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n672), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n591), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n549), .A2(KEYINPUT107), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n585), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n213), .ZN(G1324gat));
  NAND3_X1  g502(.A1(new_n591), .A2(new_n533), .A3(new_n696), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT42), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(G8gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT108), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1325gat));
  INV_X1    g510(.A(new_n373), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n697), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n362), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n697), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n697), .A2(new_n573), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  OR2_X1    g518(.A1(new_n571), .A2(new_n572), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT109), .A3(new_n587), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n573), .B2(new_n565), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n562), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n580), .A2(new_n725), .A3(new_n589), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n580), .B2(new_n589), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT44), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(KEYINPUT44), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n574), .B2(new_n590), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n627), .A2(new_n695), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n273), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n701), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n729), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n701), .A2(new_n739), .A3(G29gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n591), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(G1328gat));
  OAI21_X1  g542(.A(G36gat), .B1(new_n737), .B2(new_n586), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n739), .A2(G36gat), .A3(new_n586), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n591), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1329gat));
  INV_X1    g547(.A(new_n739), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n591), .A2(new_n227), .A3(new_n362), .A4(new_n749), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n730), .A2(new_n712), .A3(new_n732), .A4(new_n735), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n227), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT47), .B(new_n750), .C1(new_n751), .C2(new_n227), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  NOR3_X1   g555(.A1(new_n739), .A2(new_n573), .A3(G50gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n591), .A2(new_n757), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n730), .A2(new_n578), .A3(new_n732), .A4(new_n735), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT48), .B(new_n758), .C1(new_n759), .C2(new_n228), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n733), .A2(new_n720), .A3(new_n736), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n761), .A2(G50gat), .B1(new_n591), .B2(new_n757), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n762), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g562(.A(new_n695), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n672), .A2(new_n273), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n728), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n701), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g569(.A(new_n586), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n774), .A2(new_n775), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n775), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1333gat));
  OAI21_X1  g579(.A(G71gat), .B1(new_n766), .B2(new_n712), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n714), .A2(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n720), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n627), .A2(new_n273), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n728), .A2(new_n729), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT51), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n728), .A2(new_n790), .A3(new_n729), .A4(new_n787), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n695), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n632), .A2(new_n634), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n768), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n733), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n787), .A2(new_n695), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n795), .A2(new_n701), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n797), .B2(new_n793), .ZN(G1336gat));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n586), .A2(G92gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n789), .A2(new_n695), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n730), .A2(new_n586), .A3(new_n732), .A4(new_n796), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n633), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI221_X1 g605(.A(new_n801), .B1(new_n802), .B2(new_n799), .C1(new_n804), .C2(new_n633), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1337gat));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n362), .ZN(new_n809));
  INV_X1    g608(.A(G99gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n796), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n712), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(G1338gat));
  NOR2_X1   g612(.A1(new_n578), .A2(G106gat), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n789), .A2(new_n695), .A3(new_n791), .A4(new_n814), .ZN(new_n815));
  NOR4_X1   g614(.A1(new_n730), .A2(new_n573), .A3(new_n732), .A4(new_n796), .ZN(new_n816));
  INV_X1    g615(.A(G106gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NOR4_X1   g619(.A1(new_n730), .A2(new_n578), .A3(new_n732), .A4(new_n796), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n815), .B(new_n820), .C1(new_n821), .C2(new_n817), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(G1339gat));
  NOR3_X1   g622(.A1(new_n672), .A2(new_n273), .A3(new_n695), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n680), .A2(new_n686), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT10), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n646), .A2(new_n613), .A3(KEYINPUT10), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n674), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n688), .A3(KEYINPUT54), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n675), .C1(new_n679), .C2(new_n687), .ZN(new_n832));
  INV_X1    g631(.A(new_n694), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n690), .A2(new_n694), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT55), .A4(new_n833), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n269), .B2(new_n272), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n258), .A2(new_n242), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n241), .A2(new_n244), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT113), .B(new_n207), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n207), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n272), .A2(new_n695), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n671), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n839), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n846), .A2(new_n843), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n729), .A4(new_n272), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n627), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n824), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n701), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n576), .A2(new_n579), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n533), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n273), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n768), .A2(new_n586), .A3(new_n362), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n854), .B2(new_n720), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n627), .B1(new_n848), .B2(new_n851), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n862), .B(new_n573), .C1(new_n863), .C2(new_n824), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n860), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n273), .A2(G113gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n858), .B2(new_n695), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n695), .A2(G120gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n865), .B2(new_n869), .ZN(G1341gat));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  INV_X1    g670(.A(new_n865), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n853), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n281), .ZN(new_n874));
  INV_X1    g673(.A(new_n858), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n853), .A2(G127gat), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n871), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  OAI221_X1 g678(.A(KEYINPUT115), .B1(new_n875), .B2(new_n877), .C1(new_n873), .C2(new_n281), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1342gat));
  NOR2_X1   g680(.A1(new_n671), .A2(new_n533), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT116), .ZN(new_n883));
  AND4_X1   g682(.A1(new_n284), .A2(new_n855), .A3(new_n856), .A4(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n872), .B2(new_n671), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1343gat));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n273), .A2(new_n849), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n272), .A2(new_n695), .A3(new_n843), .A4(new_n846), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n729), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n851), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n853), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n824), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n578), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n888), .B1(new_n895), .B2(KEYINPUT57), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  OAI211_X1 g696(.A(KEYINPUT118), .B(new_n897), .C1(new_n854), .C2(new_n578), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n894), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT57), .A3(new_n720), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n768), .A2(new_n586), .A3(new_n712), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT117), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n273), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G141gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n712), .A2(new_n463), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT119), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n855), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n908), .A2(new_n403), .A3(new_n586), .A4(new_n273), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n903), .A2(new_n695), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT57), .B1(new_n854), .B2(new_n578), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n897), .A3(new_n720), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G148gat), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT59), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n695), .A3(new_n903), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n404), .A2(KEYINPUT59), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n908), .A2(new_n404), .A3(new_n586), .A4(new_n695), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1345gat));
  NAND3_X1  g727(.A1(new_n901), .A2(new_n627), .A3(new_n903), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G155gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n908), .A2(new_n586), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n853), .A2(G155gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1346gat));
  INV_X1    g732(.A(G162gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n901), .A2(new_n729), .A3(new_n903), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n908), .A2(new_n934), .A3(new_n883), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n854), .A2(new_n768), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n856), .A2(new_n533), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G169gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n273), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT122), .Z(new_n946));
  NAND3_X1  g745(.A1(new_n701), .A2(new_n533), .A3(new_n362), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n861), .B2(new_n864), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n948), .B2(new_n273), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n950), .A3(new_n951), .ZN(G1348gat));
  INV_X1    g751(.A(G176gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n943), .A2(new_n953), .A3(new_n695), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n948), .A2(new_n695), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n953), .ZN(G1349gat));
  AOI21_X1  g755(.A(new_n319), .B1(new_n948), .B2(new_n627), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n627), .A2(new_n288), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT125), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  INV_X1    g762(.A(new_n959), .ZN(new_n964));
  AOI211_X1 g763(.A(new_n853), .B(new_n947), .C1(new_n861), .C2(new_n864), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n963), .B(new_n964), .C1(new_n965), .C2(new_n319), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n960), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n962), .B1(new_n960), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n289), .A3(new_n729), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n948), .A2(new_n729), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(G190gat), .ZN(new_n973));
  AOI211_X1 g772(.A(KEYINPUT61), .B(new_n289), .C1(new_n948), .C2(new_n729), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n906), .A2(new_n586), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n941), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n273), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n768), .A2(new_n586), .A3(new_n373), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n916), .A2(new_n917), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n274), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n979), .A2(new_n983), .ZN(G1352gat));
  AND4_X1   g783(.A1(new_n693), .A2(new_n941), .A3(new_n695), .A4(new_n976), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  OAI21_X1  g785(.A(G204gat), .B1(new_n981), .B2(new_n764), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n978), .A2(new_n387), .A3(new_n627), .ZN(new_n993));
  OAI21_X1  g792(.A(G211gat), .B1(new_n981), .B2(new_n853), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  AOI21_X1  g797(.A(G218gat), .B1(new_n978), .B2(new_n729), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n981), .A2(new_n388), .A3(new_n671), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n999), .A2(new_n1000), .ZN(G1355gat));
endmodule


