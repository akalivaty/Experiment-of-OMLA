

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U326 ( .A(n389), .B(n294), .ZN(n391) );
  NOR2_X1 U327 ( .A1(n484), .A2(n475), .ZN(n476) );
  XNOR2_X1 U328 ( .A(n346), .B(n345), .ZN(n572) );
  XNOR2_X1 U329 ( .A(n342), .B(n341), .ZN(n344) );
  AND2_X1 U330 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U331 ( .A(G29GAT), .B(KEYINPUT71), .Z(n295) );
  NOR2_X1 U332 ( .A1(n591), .A2(n460), .ZN(n461) );
  XNOR2_X1 U333 ( .A(n391), .B(n423), .ZN(n392) );
  INV_X1 U334 ( .A(KEYINPUT90), .ZN(n398) );
  XNOR2_X1 U335 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U336 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U337 ( .A(n337), .B(n300), .ZN(n302) );
  XNOR2_X1 U338 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U339 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U340 ( .A1(n478), .A2(n450), .ZN(n451) );
  XNOR2_X1 U341 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U342 ( .A(n308), .B(n307), .ZN(n312) );
  XNOR2_X1 U343 ( .A(n488), .B(KEYINPUT120), .ZN(n583) );
  INV_X1 U344 ( .A(G43GAT), .ZN(n453) );
  XNOR2_X1 U345 ( .A(n452), .B(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U346 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U347 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U348 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U349 ( .A(n482), .B(n481), .ZN(G1355GAT) );
  XNOR2_X1 U350 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(G92GAT), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G85GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n337) );
  NAND2_X1 U355 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  INV_X1 U356 ( .A(KEYINPUT33), .ZN(n298) );
  INV_X1 U357 ( .A(KEYINPUT75), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n308) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G204GAT), .Z(n385) );
  XNOR2_X1 U360 ( .A(G120GAT), .B(n385), .ZN(n306) );
  XOR2_X1 U361 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n304) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U364 ( .A(G64GAT), .B(G78GAT), .Z(n310) );
  XNOR2_X1 U365 ( .A(G71GAT), .B(G57GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U367 ( .A(KEYINPUT13), .B(n311), .Z(n350) );
  XNOR2_X1 U368 ( .A(n312), .B(n350), .ZN(n591) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G22GAT), .Z(n314) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(G113GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U372 ( .A(G8GAT), .B(G197GAT), .Z(n316) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U375 ( .A(n318), .B(n317), .Z(n324) );
  XOR2_X1 U376 ( .A(G36GAT), .B(G43GAT), .Z(n321) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n295), .B(n319), .ZN(n336) );
  XNOR2_X1 U379 ( .A(n336), .B(G1GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U381 ( .A(G50GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n326) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT73), .Z(n330) );
  XNOR2_X1 U388 ( .A(KEYINPUT70), .B(KEYINPUT72), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n331), .B(KEYINPUT68), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n588) );
  INV_X1 U392 ( .A(n588), .ZN(n575) );
  NOR2_X1 U393 ( .A1(n591), .A2(n575), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n334), .B(KEYINPUT76), .ZN(n499) );
  XNOR2_X1 U395 ( .A(G43GAT), .B(G190GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n335), .B(G134GAT), .ZN(n378) );
  XOR2_X1 U397 ( .A(n336), .B(n378), .Z(n338) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U399 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n342) );
  NAND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  INV_X1 U401 ( .A(KEYINPUT9), .ZN(n339) );
  XOR2_X1 U402 ( .A(G36GAT), .B(G218GAT), .Z(n431) );
  XOR2_X1 U403 ( .A(G50GAT), .B(G162GAT), .Z(n389) );
  XNOR2_X1 U404 ( .A(n431), .B(n389), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n572), .B(KEYINPUT77), .ZN(n489) );
  XNOR2_X1 U407 ( .A(KEYINPUT36), .B(n489), .ZN(n478) );
  XOR2_X1 U408 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n348) );
  XOR2_X1 U409 ( .A(G15GAT), .B(G127GAT), .Z(n365) );
  XOR2_X1 U410 ( .A(G8GAT), .B(G211GAT), .Z(n430) );
  XNOR2_X1 U411 ( .A(n365), .B(n430), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U413 ( .A(n349), .B(KEYINPUT81), .Z(n352) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U416 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n354) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U419 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n358) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(KEYINPUT12), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G155GAT), .Z(n386) );
  XNOR2_X1 U424 ( .A(n359), .B(n386), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n568) );
  XOR2_X1 U426 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n363) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G71GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U429 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U430 ( .A1(G227GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n369) );
  XNOR2_X1 U433 ( .A(KEYINPUT65), .B(KEYINPUT87), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n372) );
  XOR2_X1 U435 ( .A(G120GAT), .B(KEYINPUT83), .Z(n371) );
  XNOR2_X1 U436 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n407) );
  XOR2_X1 U438 ( .A(n372), .B(n407), .Z(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n374) );
  XNOR2_X1 U440 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U442 ( .A(n375), .B(G176GAT), .Z(n377) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n435) );
  XNOR2_X1 U445 ( .A(n435), .B(n378), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U447 ( .A(n382), .B(n381), .Z(n543) );
  XNOR2_X1 U448 ( .A(n543), .B(KEYINPUT89), .ZN(n437) );
  XOR2_X1 U449 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n384) );
  XNOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n403) );
  XOR2_X1 U452 ( .A(n385), .B(G211GAT), .Z(n388) );
  XNOR2_X1 U453 ( .A(G78GAT), .B(n386), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n393) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n390), .B(KEYINPUT91), .ZN(n423) );
  XOR2_X1 U457 ( .A(n393), .B(n392), .Z(n395) );
  XNOR2_X1 U458 ( .A(G218GAT), .B(G106GAT), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n401) );
  XOR2_X1 U460 ( .A(KEYINPUT92), .B(KEYINPUT3), .Z(n397) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n406), .B(KEYINPUT22), .ZN(n399) );
  XOR2_X1 U464 ( .A(n403), .B(n402), .Z(n483) );
  XNOR2_X1 U465 ( .A(n483), .B(KEYINPUT28), .ZN(n546) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT96), .B(KEYINPUT4), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n422) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n420) );
  XOR2_X1 U470 ( .A(G85GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U471 ( .A(G29GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U473 ( .A(G148GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G127GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U476 ( .A(n413), .B(n412), .Z(n418) );
  XOR2_X1 U477 ( .A(KEYINPUT5), .B(G57GAT), .Z(n415) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U480 ( .A(KEYINPUT95), .B(n416), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n517) );
  INV_X1 U484 ( .A(n517), .ZN(n532) );
  XOR2_X1 U485 ( .A(KEYINPUT97), .B(n423), .Z(n425) );
  NAND2_X1 U486 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U488 ( .A(G204GAT), .B(G64GAT), .Z(n427) );
  XNOR2_X1 U489 ( .A(G190GAT), .B(G92GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U491 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n534) );
  XOR2_X1 U495 ( .A(KEYINPUT27), .B(n534), .Z(n440) );
  NAND2_X1 U496 ( .A1(n532), .A2(n440), .ZN(n541) );
  NOR2_X1 U497 ( .A1(n546), .A2(n541), .ZN(n436) );
  NAND2_X1 U498 ( .A1(n437), .A2(n436), .ZN(n449) );
  INV_X1 U499 ( .A(n543), .ZN(n523) );
  NAND2_X1 U500 ( .A1(n483), .A2(n523), .ZN(n439) );
  XNOR2_X1 U501 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n475) );
  INV_X1 U503 ( .A(n475), .ZN(n562) );
  NAND2_X1 U504 ( .A1(n562), .A2(n440), .ZN(n441) );
  XOR2_X1 U505 ( .A(KEYINPUT99), .B(n441), .Z(n446) );
  NOR2_X1 U506 ( .A1(n534), .A2(n523), .ZN(n442) );
  NOR2_X1 U507 ( .A1(n483), .A2(n442), .ZN(n443) );
  XNOR2_X1 U508 ( .A(KEYINPUT25), .B(n443), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n444), .B(KEYINPUT100), .ZN(n445) );
  NAND2_X1 U510 ( .A1(n446), .A2(n445), .ZN(n447) );
  NAND2_X1 U511 ( .A1(n447), .A2(n517), .ZN(n448) );
  NAND2_X1 U512 ( .A1(n449), .A2(n448), .ZN(n497) );
  NAND2_X1 U513 ( .A1(n568), .A2(n497), .ZN(n450) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n451), .Z(n529) );
  NAND2_X1 U515 ( .A1(n499), .A2(n529), .ZN(n452) );
  NOR2_X1 U516 ( .A1(n514), .A2(n523), .ZN(n456) );
  XNOR2_X1 U517 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n454) );
  NOR2_X1 U518 ( .A1(n568), .A2(n478), .ZN(n458) );
  XNOR2_X1 U519 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U521 ( .A(n459), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT111), .ZN(n462) );
  NOR2_X1 U523 ( .A1(n462), .A2(n588), .ZN(n463) );
  XNOR2_X1 U524 ( .A(KEYINPUT112), .B(n463), .ZN(n470) );
  INV_X1 U525 ( .A(KEYINPUT41), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(n591), .ZN(n549) );
  NAND2_X1 U527 ( .A1(n549), .A2(n588), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT46), .ZN(n466) );
  XNOR2_X1 U529 ( .A(KEYINPUT110), .B(n568), .ZN(n582) );
  NAND2_X1 U530 ( .A1(n466), .A2(n582), .ZN(n467) );
  NOR2_X1 U531 ( .A1(n572), .A2(n467), .ZN(n468) );
  XOR2_X1 U532 ( .A(KEYINPUT47), .B(n468), .Z(n469) );
  NOR2_X1 U533 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U535 ( .A1(n542), .A2(n534), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n472), .B(KEYINPUT54), .ZN(n473) );
  NAND2_X1 U537 ( .A1(n473), .A2(n517), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n474), .B(KEYINPUT64), .ZN(n484) );
  XOR2_X1 U539 ( .A(n476), .B(KEYINPUT123), .Z(n595) );
  INV_X1 U540 ( .A(n595), .ZN(n477) );
  NOR2_X1 U541 ( .A1(n478), .A2(n477), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n480) );
  INV_X1 U543 ( .A(G218GAT), .ZN(n479) );
  NOR2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  NAND2_X1 U547 ( .A1(n487), .A2(n543), .ZN(n488) );
  INV_X1 U548 ( .A(n489), .ZN(n490) );
  INV_X1 U549 ( .A(n490), .ZN(n556) );
  NOR2_X1 U550 ( .A1(n583), .A2(n556), .ZN(n494) );
  XNOR2_X1 U551 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n492) );
  INV_X1 U552 ( .A(G190GAT), .ZN(n491) );
  INV_X1 U553 ( .A(n568), .ZN(n594) );
  NAND2_X1 U554 ( .A1(n594), .A2(n556), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(n495), .Z(n496) );
  NAND2_X1 U556 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(KEYINPUT101), .ZN(n516) );
  NAND2_X1 U558 ( .A1(n516), .A2(n499), .ZN(n506) );
  NOR2_X1 U559 ( .A1(n517), .A2(n506), .ZN(n500) );
  XOR2_X1 U560 ( .A(G1GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U561 ( .A(KEYINPUT34), .B(n501), .ZN(G1324GAT) );
  NOR2_X1 U562 ( .A1(n534), .A2(n506), .ZN(n502) );
  XOR2_X1 U563 ( .A(G8GAT), .B(n502), .Z(G1325GAT) );
  NOR2_X1 U564 ( .A1(n523), .A2(n506), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(n505), .ZN(G1326GAT) );
  INV_X1 U568 ( .A(n546), .ZN(n526) );
  NOR2_X1 U569 ( .A1(n526), .A2(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G22GAT), .B(n509), .ZN(G1327GAT) );
  NOR2_X1 U573 ( .A1(n514), .A2(n517), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G29GAT), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n514), .A2(n534), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1329GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n514), .ZN(n515) );
  XOR2_X1 U580 ( .A(G50GAT), .B(n515), .Z(G1331GAT) );
  INV_X1 U581 ( .A(n549), .ZN(n577) );
  NOR2_X1 U582 ( .A1(n588), .A2(n577), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n530), .A2(n516), .ZN(n525) );
  NOR2_X1 U584 ( .A1(n517), .A2(n525), .ZN(n519) );
  XNOR2_X1 U585 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G57GAT), .B(n520), .ZN(G1332GAT) );
  NOR2_X1 U588 ( .A1(n534), .A2(n525), .ZN(n521) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(n521), .Z(n522) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(n522), .ZN(G1333GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n525), .ZN(n524) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n524), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT109), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n532), .A2(n538), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n533), .ZN(G1336GAT) );
  INV_X1 U600 ( .A(n534), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n535), .A2(n538), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G92GAT), .B(n536), .ZN(G1337GAT) );
  NAND2_X1 U603 ( .A1(n538), .A2(n543), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n561) );
  NAND2_X1 U609 ( .A1(n543), .A2(n561), .ZN(n544) );
  XOR2_X1 U610 ( .A(KEYINPUT113), .B(n544), .Z(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT114), .B(n547), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n588), .A2(n552), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(n548), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n552), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  INV_X1 U618 ( .A(n552), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n555), .A2(n582), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT50), .B(n553), .Z(n554) );
  XNOR2_X1 U621 ( .A(G127GAT), .B(n554), .ZN(G1342GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n558) );
  XNOR2_X1 U624 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1343GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n571) );
  NOR2_X1 U628 ( .A1(n575), .A2(n571), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1344GAT) );
  NOR2_X1 U631 ( .A1(n577), .A2(n571), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G148GAT), .B(n567), .ZN(G1345GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n571), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT118), .B(n569), .Z(n570) );
  XNOR2_X1 U637 ( .A(G155GAT), .B(n570), .ZN(G1346GAT) );
  INV_X1 U638 ( .A(n571), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n576) );
  XOR2_X1 U642 ( .A(G169GAT), .B(n576), .Z(G1348GAT) );
  NOR2_X1 U643 ( .A1(n577), .A2(n583), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n579) );
  XNOR2_X1 U645 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1349GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G183GAT), .B(n584), .Z(G1350GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT60), .B(n587), .Z(n590) );
  NAND2_X1 U654 ( .A1(n595), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  XOR2_X1 U656 ( .A(G204GAT), .B(KEYINPUT61), .Z(n593) );
  NAND2_X1 U657 ( .A1(n595), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G211GAT), .B(n596), .ZN(G1354GAT) );
endmodule

