//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G116), .A2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n217), .B(new_n222), .C1(G97), .C2(G257), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n211), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(new_n203), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n248), .B1(new_n249), .B2(new_n251), .C1(new_n252), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n226), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n202), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n262), .A2(new_n258), .A3(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G20), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT68), .B1(new_n262), .B2(new_n258), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(new_n202), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(G222), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n253), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n280), .B(new_n283), .C1(G77), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n282), .A2(new_n286), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n285), .B(new_n289), .C1(new_n219), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n269), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(new_n295), .B1(G200), .B2(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n272), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n272), .A2(new_n299), .A3(new_n293), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n291), .A2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n294), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  INV_X1    g0106(.A(G232), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G226), .B2(G1698), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n306), .B1(new_n309), .B2(new_n276), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n283), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n282), .A2(G238), .A3(new_n286), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n289), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(new_n303), .B1(KEYINPUT71), .B2(KEYINPUT14), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n319));
  INV_X1    g0119(.A(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n314), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(G169), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(G179), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n318), .A2(new_n319), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n220), .A2(G20), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n326), .B1(new_n251), .B2(new_n202), .C1(new_n255), .C2(new_n213), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT70), .B(KEYINPUT11), .Z(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n258), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n327), .B2(new_n258), .ZN(new_n330));
  INV_X1    g0130(.A(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(G13), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G1), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n258), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G68), .A3(new_n265), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT12), .B1(new_n331), .B2(new_n333), .ZN(new_n338));
  NOR4_X1   g0138(.A1(new_n329), .A2(new_n330), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n325), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n317), .B2(G190), .ZN(new_n342));
  INV_X1    g0142(.A(G200), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n317), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n276), .B1(G232), .B2(new_n277), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n221), .B2(new_n277), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n283), .C1(G107), .C2(new_n284), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n289), .C1(new_n214), .C2(new_n290), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(G179), .ZN(new_n350));
  INV_X1    g0150(.A(new_n252), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT15), .B(G87), .Z(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n250), .B1(new_n352), .B2(new_n254), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n208), .B2(new_n213), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n258), .B1(new_n213), .B2(new_n262), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n335), .A2(G77), .A3(new_n265), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n349), .A2(new_n303), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n345), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n301), .A2(new_n305), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n250), .A2(G159), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G58), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n220), .ZN(new_n368));
  OAI21_X1  g0168(.A(G20), .B1(new_n368), .B2(new_n201), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n284), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n220), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n363), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n370), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT72), .B1(new_n274), .B2(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n275), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n274), .A2(KEYINPUT72), .A3(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n208), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n381), .B2(KEYINPUT7), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n380), .B2(new_n208), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n376), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n375), .B(new_n258), .C1(new_n384), .C2(new_n363), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n290), .A2(new_n307), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n274), .A2(KEYINPUT72), .A3(G33), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n275), .B2(new_n377), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n219), .A2(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n279), .A2(new_n277), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI211_X1 g0193(.A(new_n386), .B(new_n288), .C1(new_n393), .C2(new_n283), .ZN(new_n394));
  XOR2_X1   g0194(.A(KEYINPUT74), .B(G190), .Z(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n283), .ZN(new_n397));
  INV_X1    g0197(.A(new_n386), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n289), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G200), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n351), .A2(new_n261), .ZN(new_n401));
  INV_X1    g0201(.A(new_n267), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n351), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n385), .A2(new_n396), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n385), .A2(new_n403), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n397), .A2(G179), .A3(new_n398), .A4(new_n289), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n394), .B2(new_n303), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(KEYINPUT18), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n349), .A2(G200), .ZN(new_n414));
  INV_X1    g0214(.A(new_n357), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n292), .C2(new_n349), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n362), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n207), .A2(G33), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n335), .A2(KEYINPUT75), .A3(new_n261), .A4(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n261), .A2(new_n420), .A3(new_n226), .A4(new_n257), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n424), .A3(G107), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n333), .A2(G20), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT25), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(KEYINPUT25), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT81), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n425), .A2(new_n432), .A3(new_n428), .A4(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n215), .A2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n284), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT22), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT23), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n208), .B2(G107), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n426), .A2(KEYINPUT23), .A3(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n436), .A2(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n254), .A2(G116), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT22), .A4(new_n435), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n441), .A2(KEYINPUT24), .A3(new_n442), .A4(new_n443), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n258), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n434), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G45), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(G264), .A3(new_n282), .ZN(new_n455));
  INV_X1    g0255(.A(G257), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n216), .A2(new_n277), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n378), .A2(new_n379), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n455), .B1(new_n461), .B2(new_n283), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n451), .B(G274), .C1(new_n453), .C2(new_n452), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n303), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G179), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n449), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n462), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT82), .B1(new_n462), .B2(new_n464), .ZN(new_n475));
  OAI21_X1  g0275(.A(G169), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n471), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(new_n434), .B2(new_n448), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n208), .B1(new_n483), .B2(G33), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT78), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT78), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT79), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n208), .A2(G116), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n226), .B2(new_n257), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n422), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n333), .B2(new_n494), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n487), .A2(new_n495), .A3(new_n490), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT79), .A2(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n492), .A2(new_n493), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n277), .A2(G264), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n456), .A2(new_n277), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n378), .A2(new_n379), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n276), .A2(G303), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n454), .A2(G270), .A3(new_n282), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n464), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n504), .A2(new_n512), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(G200), .ZN(new_n516));
  INV_X1    g0316(.A(new_n504), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n395), .A3(new_n464), .A4(new_n511), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n512), .A2(new_n470), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n504), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n504), .A2(new_n512), .A3(KEYINPUT21), .A4(G169), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n515), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT80), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n343), .A2(KEYINPUT77), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n273), .A2(new_n275), .A3(G250), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n277), .B1(new_n527), .B2(KEYINPUT4), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n276), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n528), .A2(new_n486), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n380), .B2(new_n214), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n282), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n454), .A2(new_n282), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n464), .B1(new_n456), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n526), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n421), .A2(new_n424), .A3(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n483), .A2(new_n426), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n426), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n208), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n251), .A2(new_n213), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n372), .A2(new_n373), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n548), .C1(new_n549), .C2(new_n426), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n539), .B1(new_n550), .B2(new_n258), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n262), .A2(new_n483), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n532), .B1(new_n284), .B2(G250), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n485), .B(new_n553), .C1(new_n554), .C2(new_n277), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT4), .B1(new_n388), .B2(G244), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n283), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n535), .A2(new_n456), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT77), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n292), .B1(new_n562), .B2(new_n343), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n537), .A2(new_n551), .A3(new_n552), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n303), .B1(new_n534), .B2(new_n536), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n426), .B1(new_n372), .B2(new_n373), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n567), .A2(new_n547), .A3(new_n545), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n552), .B(new_n538), .C1(new_n568), .C2(new_n335), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n557), .A2(new_n561), .A3(new_n470), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n434), .A2(new_n448), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n474), .A2(new_n475), .A3(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n465), .A2(new_n343), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n214), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n221), .A2(new_n277), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n378), .A2(new_n379), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G116), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n283), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n207), .A2(G45), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n282), .A2(G250), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n287), .B2(new_n584), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n587), .A3(G190), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n282), .B1(new_n580), .B2(new_n581), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n589), .B2(new_n586), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n378), .A2(new_n379), .A3(new_n208), .A4(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n208), .A3(G33), .A4(G97), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G87), .A2(G97), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n426), .B1(new_n306), .B2(new_n208), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n352), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n258), .B1(new_n262), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n421), .A2(new_n424), .A3(G87), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n588), .A2(new_n590), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n258), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n262), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n421), .A2(new_n424), .A3(new_n352), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n583), .A2(new_n587), .A3(new_n470), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n303), .B1(new_n589), .B2(new_n586), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n572), .A2(new_n577), .A3(new_n609), .ZN(new_n610));
  NOR4_X1   g0410(.A1(new_n419), .A2(new_n482), .A3(new_n525), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n305), .ZN(new_n612));
  INV_X1    g0412(.A(new_n413), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n360), .A2(new_n344), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n341), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n405), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n612), .B1(new_n617), .B2(new_n301), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n515), .A2(new_n521), .A3(new_n522), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n478), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n610), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n609), .A2(new_n571), .A3(new_n565), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n467), .A2(new_n292), .A3(new_n468), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n449), .B1(new_n625), .B2(new_n575), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n620), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n472), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT84), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n609), .A3(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n601), .A2(new_n608), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n571), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(new_n608), .ZN(new_n638));
  INV_X1    g0438(.A(new_n608), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT85), .B(new_n639), .C1(new_n633), .C2(new_n636), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n623), .A2(new_n630), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n619), .B1(new_n418), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT86), .ZN(G369));
  NOR2_X1   g0443(.A1(new_n482), .A2(new_n626), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n332), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n207), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G343), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n628), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n650), .B(KEYINPUT89), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n644), .A2(new_n652), .B1(new_n478), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n504), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n523), .B(KEYINPUT80), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n656), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT87), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n644), .B1(new_n573), .B2(new_n650), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n472), .B2(new_n650), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n662), .B2(new_n665), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n655), .B1(new_n667), .B2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n209), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n594), .A2(new_n426), .A3(new_n497), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n672), .A3(new_n207), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n229), .B2(new_n671), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  INV_X1    g0475(.A(KEYINPUT29), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n608), .B(KEYINPUT91), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n620), .B1(new_n473), .B2(new_n480), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n637), .B(new_n677), .C1(new_n678), .C2(new_n610), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n676), .B1(new_n679), .B2(new_n650), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT26), .B1(new_n632), .B2(new_n609), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n571), .A2(new_n635), .A3(new_n634), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n608), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT85), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n637), .A2(new_n631), .A3(new_n608), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n622), .B1(new_n610), .B2(new_n621), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n627), .A2(new_n629), .A3(KEYINPUT84), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n681), .B1(new_n689), .B2(new_n653), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n641), .A2(KEYINPUT90), .A3(new_n654), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n680), .B1(new_n692), .B2(new_n676), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n658), .A2(new_n481), .A3(new_n627), .A4(new_n654), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n534), .A2(new_n536), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n589), .A2(new_n586), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n520), .A2(new_n696), .A3(new_n462), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n557), .A2(new_n561), .ZN(new_n702));
  AND4_X1   g0502(.A1(new_n470), .A2(new_n702), .A3(new_n465), .A4(new_n512), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n583), .A2(new_n587), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n699), .A2(new_n700), .B1(new_n704), .B2(new_n703), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n650), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n695), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n694), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n675), .B1(new_n714), .B2(G1), .ZN(G364));
  INV_X1    g0515(.A(new_n671), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n645), .A2(G45), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n662), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n660), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(G20), .A3(new_n292), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n284), .B1(new_n724), .B2(G329), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n208), .A2(new_n470), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n727), .A2(new_n343), .A3(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT33), .B(G317), .Z(new_n730));
  OAI21_X1  g0530(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n395), .A2(new_n726), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n343), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(G326), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G311), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n208), .A2(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(G303), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n208), .B1(new_n722), .B2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(G294), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n737), .A2(new_n292), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(G283), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n732), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G322), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n734), .A2(new_n736), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n740), .A2(new_n483), .ZN(new_n749));
  INV_X1    g0549(.A(new_n735), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n284), .B1(new_n750), .B2(new_n213), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n749), .B(new_n751), .C1(G107), .C2(new_n744), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G50), .A2(new_n733), .B1(new_n746), .B2(G58), .ZN(new_n753));
  INV_X1    g0553(.A(new_n738), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G87), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n723), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n757), .B(new_n758), .Z(new_n759));
  NAND4_X1  g0559(.A1(new_n752), .A2(new_n753), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n729), .A2(new_n220), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n748), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n226), .B1(G20), .B2(new_n303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT92), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n763), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n388), .A2(new_n670), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n229), .A2(new_n450), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n243), .C2(new_n450), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n284), .A2(new_n209), .A3(G355), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(G116), .C2(new_n209), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n762), .A2(new_n763), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n767), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n719), .B(new_n774), .C1(new_n660), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n721), .A2(new_n776), .ZN(G396));
  OAI21_X1  g0577(.A(new_n416), .B1(new_n415), .B2(new_n650), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n359), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n360), .A2(new_n650), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n641), .A2(new_n654), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n692), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(new_n713), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n718), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n388), .B1(new_n367), .B2(new_n740), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n744), .A2(G68), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n202), .B2(new_n738), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT94), .Z(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n746), .A2(G143), .B1(G150), .B2(new_n728), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  INV_X1    g0593(.A(new_n733), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n793), .B2(new_n794), .C1(new_n756), .C2(new_n750), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n787), .B(new_n790), .C1(new_n791), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n791), .B2(new_n795), .C1(new_n797), .C2(new_n723), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n723), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n276), .B1(new_n750), .B2(new_n497), .C1(new_n801), .C2(new_n729), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G303), .B2(new_n733), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n743), .A2(new_n215), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n749), .B(new_n804), .C1(G107), .C2(new_n754), .ZN(new_n805));
  INV_X1    g0605(.A(new_n746), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n803), .B(new_n805), .C1(new_n741), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n798), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n763), .A2(new_n764), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n808), .A2(new_n763), .B1(new_n213), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n810), .B(new_n719), .C1(new_n782), .C2(new_n766), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n786), .A2(new_n811), .ZN(G384));
  AOI21_X1  g0612(.A(new_n619), .B1(new_n694), .B2(new_n418), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n405), .A2(new_n413), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT97), .ZN(new_n815));
  INV_X1    g0615(.A(new_n403), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n388), .A2(G20), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n220), .B1(new_n817), .B2(new_n371), .ZN(new_n818));
  INV_X1    g0618(.A(new_n383), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n370), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n335), .B1(new_n820), .B2(KEYINPUT16), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n384), .A2(new_n363), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n649), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n815), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n822), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n258), .B1(new_n384), .B2(new_n363), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n403), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(KEYINPUT97), .A3(new_n649), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n814), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(new_n408), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n825), .A2(new_n829), .A3(new_n404), .A4(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n406), .B1(new_n408), .B2(new_n649), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n404), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(KEYINPUT37), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n831), .B(KEYINPUT38), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n833), .B2(KEYINPUT37), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n405), .A2(new_n413), .B1(new_n825), .B2(new_n829), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n345), .A2(new_n340), .A3(new_n651), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n341), .B(new_n344), .C1(new_n339), .C2(new_n650), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n783), .A2(KEYINPUT96), .A3(new_n780), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT96), .B1(new_n783), .B2(new_n780), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n844), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n836), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n406), .A2(new_n649), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n405), .B2(new_n413), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n839), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT39), .B1(new_n838), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n341), .A2(new_n651), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n851), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n613), .A2(new_n824), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n850), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n813), .B(new_n862), .Z(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n695), .A2(new_n710), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n847), .A3(new_n782), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n843), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n866), .A2(new_n847), .A3(new_n782), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n838), .A2(new_n856), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n418), .A2(new_n866), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G330), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n863), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n207), .B2(new_n645), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n543), .A2(new_n544), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT95), .Z(new_n880));
  AOI21_X1  g0680(.A(new_n497), .B1(new_n880), .B2(KEYINPUT35), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(new_n227), .C1(KEYINPUT35), .C2(new_n880), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT36), .ZN(new_n883));
  OAI21_X1  g0683(.A(G77), .B1(new_n367), .B2(new_n220), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n884), .A2(new_n228), .B1(G50), .B2(new_n220), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(G1), .A3(new_n332), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n878), .A2(new_n883), .A3(new_n886), .ZN(G367));
  INV_X1    g0687(.A(new_n668), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n653), .A2(new_n569), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n572), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n571), .B2(new_n654), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT99), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n888), .A2(new_n666), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n644), .A2(new_n652), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT42), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n632), .B1(new_n893), .B2(new_n482), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n897), .B1(new_n653), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT43), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n650), .B1(new_n599), .B2(new_n600), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n608), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n609), .B2(new_n901), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT98), .Z(new_n904));
  OAI211_X1 g0704(.A(new_n894), .B(new_n899), .C1(new_n900), .C2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n904), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n899), .B1(new_n900), .B2(new_n904), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n908), .A2(new_n666), .A3(new_n888), .A4(new_n893), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(KEYINPUT43), .B2(new_n906), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n671), .B(KEYINPUT41), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n662), .A2(KEYINPUT100), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n895), .B1(new_n665), .B2(new_n652), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT100), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n661), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(KEYINPUT101), .A3(new_n714), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT101), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n918), .A2(new_n916), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n661), .B(KEYINPUT100), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  INV_X1    g0725(.A(new_n714), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n893), .A2(new_n655), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n893), .A2(new_n655), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT45), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n888), .A2(new_n929), .A3(new_n666), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n667), .B2(new_n668), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n921), .A2(new_n927), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n914), .B1(new_n937), .B2(new_n714), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n717), .A2(G1), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n910), .B(new_n912), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n738), .A2(new_n497), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n746), .A2(G303), .B1(KEYINPUT46), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n799), .B2(new_n794), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n735), .A2(G283), .B1(G317), .B2(new_n724), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(KEYINPUT46), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n729), .A2(new_n741), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n380), .B1(new_n483), .B2(new_n743), .C1(new_n426), .C2(new_n740), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n943), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G50), .A2(new_n735), .B1(new_n728), .B2(G159), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT102), .Z(new_n950));
  INV_X1    g0750(.A(G143), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n950), .B1(new_n951), .B2(new_n794), .C1(new_n249), .C2(new_n806), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n740), .A2(new_n220), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n738), .A2(new_n367), .B1(new_n793), .B2(new_n723), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(KEYINPUT103), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT103), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n744), .A2(G77), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR4_X1   g0758(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n948), .B1(new_n959), .B2(new_n284), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  AOI21_X1  g0761(.A(new_n718), .B1(new_n961), .B2(new_n763), .ZN(new_n962));
  INV_X1    g0762(.A(new_n769), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n768), .B1(new_n209), .B2(new_n598), .C1(new_n238), .C2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n962), .B(new_n964), .C1(new_n775), .C2(new_n906), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n940), .A2(new_n965), .ZN(G387));
  NAND2_X1  g0766(.A1(new_n921), .A2(new_n927), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n671), .C1(new_n714), .C2(new_n920), .ZN(new_n968));
  INV_X1    g0768(.A(new_n763), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n746), .A2(G317), .B1(G311), .B2(new_n728), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n733), .A2(G322), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(new_n739), .C2(new_n750), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT48), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n801), .B2(new_n740), .C1(new_n741), .C2(new_n738), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT49), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n724), .A2(G326), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n975), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n388), .B1(G116), .B2(new_n744), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n729), .A2(new_n252), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n735), .A2(G68), .B1(G150), .B2(new_n724), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n806), .B2(new_n202), .C1(new_n756), .C2(new_n794), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n738), .A2(new_n213), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n388), .B1(new_n483), .B2(new_n743), .C1(new_n598), .C2(new_n740), .ZN(new_n985));
  OR4_X1    g0785(.A1(new_n981), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n969), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n284), .A2(new_n209), .A3(new_n672), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n235), .A2(G45), .ZN(new_n989));
  AOI211_X1 g0789(.A(G45), .B(new_n672), .C1(G68), .C2(G77), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n252), .A2(KEYINPUT50), .A3(G50), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT50), .B1(new_n252), .B2(G50), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n769), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n988), .B1(G107), .B2(new_n209), .C1(new_n989), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n987), .B1(new_n768), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n719), .C1(new_n665), .C2(new_n775), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n920), .B2(new_n939), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n968), .A2(new_n1001), .ZN(G393));
  NAND3_X1  g0802(.A1(new_n967), .A2(new_n933), .A3(new_n935), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n671), .A3(new_n937), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n892), .A2(new_n767), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n768), .B1(new_n483), .B2(new_n209), .C1(new_n246), .C2(new_n963), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G311), .A2(new_n746), .B1(new_n733), .B2(G317), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT52), .Z(new_n1008));
  OAI22_X1  g0808(.A1(new_n729), .A2(new_n739), .B1(new_n740), .B2(new_n497), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT105), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n743), .A2(new_n426), .B1(new_n738), .B2(new_n801), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n284), .B(new_n1013), .C1(G322), .C2(new_n724), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1008), .B(new_n1015), .C1(new_n741), .C2(new_n750), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n249), .A2(new_n794), .B1(new_n806), .B2(new_n756), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT51), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n388), .B1(new_n220), .B2(new_n738), .C1(new_n215), .C2(new_n743), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n750), .A2(new_n252), .B1(new_n723), .B2(new_n951), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G50), .C2(new_n728), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n740), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(G77), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT106), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n718), .B1(new_n1028), .B2(new_n763), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1005), .A2(new_n1006), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n936), .B2(new_n939), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1004), .A2(new_n1031), .ZN(G390));
  NOR2_X1   g0832(.A1(new_n867), .A2(new_n875), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n857), .B1(new_n843), .B2(KEYINPUT39), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n859), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n679), .A2(new_n650), .A3(new_n779), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1038), .A2(new_n780), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n847), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n870), .A2(new_n1036), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1033), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n711), .A2(new_n847), .A3(G330), .A4(new_n782), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT96), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n685), .A2(new_n686), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n687), .A2(new_n688), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n653), .B(new_n781), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n780), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n783), .A2(KEYINPUT96), .A3(new_n780), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n859), .B1(new_n1054), .B2(new_n847), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1045), .B(new_n1046), .C1(new_n1055), .C2(new_n1034), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1044), .A2(new_n1056), .A3(new_n939), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n809), .A2(new_n252), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G97), .A2(new_n735), .B1(new_n728), .B2(G107), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT110), .Z(new_n1060));
  AOI22_X1  g0860(.A1(G116), .A2(new_n746), .B1(new_n733), .B2(G283), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n788), .B(new_n1024), .C1(new_n741), .C2(new_n723), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n284), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n755), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(G128), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1065), .A2(new_n794), .B1(new_n806), .B2(new_n797), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  AOI21_X1  g0867(.A(new_n276), .B1(new_n735), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n793), .B2(new_n729), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n743), .A2(new_n202), .B1(new_n740), .B2(new_n756), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n738), .A2(new_n249), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT109), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT53), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(G125), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n723), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1064), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT111), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n718), .B1(new_n1080), .B2(new_n763), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1058), .B(new_n1081), .C1(new_n1034), .C2(new_n766), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1040), .B1(new_n712), .B2(new_n781), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n875), .B2(new_n867), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n866), .A2(KEYINPUT107), .A3(G330), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n782), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT107), .B1(new_n866), .B2(G330), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1040), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1054), .A2(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n418), .A2(G330), .A3(new_n866), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n618), .B(new_n1091), .C1(new_n693), .C2(new_n419), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1044), .A2(new_n1056), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1044), .B2(new_n1056), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1097), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT108), .B1(new_n1097), .B2(new_n671), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1057), .B(new_n1082), .C1(new_n1098), .C2(new_n1099), .ZN(G378));
  NAND3_X1  g0900(.A1(new_n868), .A2(new_n871), .A3(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n862), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n850), .A3(new_n860), .A4(new_n861), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n269), .A2(new_n824), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT112), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n301), .A2(new_n1107), .A3(new_n305), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n301), .B2(new_n305), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1110), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1106), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n1108), .A3(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1105), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1103), .A2(new_n1118), .A3(new_n1104), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(KEYINPUT57), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1092), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1094), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT113), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT113), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1094), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1122), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT114), .B1(new_n1128), .B2(new_n716), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1121), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1118), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1094), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1126), .B1(new_n1094), .B2(new_n1123), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT57), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1130), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT114), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n671), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1129), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n794), .A2(new_n497), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n281), .B1(new_n723), .B2(new_n801), .C1(new_n750), .C2(new_n598), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G107), .C2(new_n746), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n743), .A2(new_n367), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n984), .A2(new_n1146), .A3(new_n388), .A4(new_n953), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n483), .C2(new_n729), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT58), .Z(new_n1149));
  OAI22_X1  g0949(.A1(new_n750), .A2(new_n793), .B1(new_n740), .B2(new_n249), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n754), .B2(new_n1067), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n1077), .B2(new_n794), .C1(new_n1065), .C2(new_n806), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G132), .B2(new_n728), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G33), .B1(new_n724), .B2(G124), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G41), .B(new_n1156), .C1(G159), .C2(new_n744), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n281), .B1(new_n380), .B2(new_n253), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1149), .B(new_n1157), .C1(new_n202), .C2(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n719), .B1(new_n969), .B2(new_n1159), .C1(new_n1118), .C2(new_n766), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n202), .B2(new_n809), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1132), .B2(new_n939), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1142), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT115), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G375));
  OAI221_X1 g0965(.A(new_n957), .B1(new_n483), .B2(new_n738), .C1(new_n598), .C2(new_n740), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n276), .B1(new_n729), .B2(new_n497), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G303), .B2(new_n724), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n801), .B2(new_n806), .C1(new_n741), .C2(new_n794), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1166), .B(new_n1169), .C1(G107), .C2(new_n735), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n380), .B(new_n1146), .C1(G50), .C2(new_n1023), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n756), .B2(new_n738), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n735), .A2(G150), .B1(G128), .B2(new_n724), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n806), .B2(new_n793), .C1(new_n797), .C2(new_n794), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(new_n728), .C2(new_n1067), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n969), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n718), .B1(new_n220), .B2(new_n809), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT117), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n1040), .C2(new_n764), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1090), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n939), .B(KEYINPUT116), .Z(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n913), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1185), .B2(new_n1093), .ZN(G381));
  NAND2_X1  g0986(.A1(new_n1057), .A2(new_n1082), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1097), .B2(new_n671), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(G375), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(G396), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n968), .A2(new_n1191), .A3(new_n1001), .ZN(new_n1192));
  OR2_X1    g0992(.A1(G381), .A2(G384), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(G387), .A2(G390), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1194), .ZN(G407));
  INV_X1    g0995(.A(G343), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1190), .B1(new_n1196), .B2(new_n1194), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(G213), .ZN(G409));
  INV_X1    g0998(.A(KEYINPUT126), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1142), .A2(G378), .A3(new_n1162), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n913), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1182), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1130), .B(new_n1131), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1188), .B1(new_n1203), .B2(new_n1161), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(G213), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(G343), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT123), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1210), .B(new_n1207), .C1(new_n1200), .C2(new_n1204), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT60), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n671), .B1(new_n1184), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT60), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1213), .A2(new_n1093), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G384), .B1(new_n1215), .B2(new_n1183), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT119), .Z(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(G384), .A3(new_n1183), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT118), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1207), .A2(G2897), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1217), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1209), .A2(new_n1211), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1199), .B1(new_n1225), .B2(KEYINPUT61), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1207), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT62), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(KEYINPUT62), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1210), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1224), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1227), .A2(KEYINPUT123), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(KEYINPUT126), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1226), .A2(new_n1233), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(new_n1192), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  AND3_X1   g1046(.A1(G387), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(G387), .B2(new_n1246), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n940), .A2(G390), .A3(new_n965), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT121), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1244), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1244), .A2(new_n1250), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G387), .B2(new_n1246), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1241), .A2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1229), .A2(KEYINPUT63), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT124), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n1257), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1239), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1230), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1262), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1256), .B1(new_n1268), .B2(new_n1269), .ZN(G405));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1200), .B1(new_n1164), .B2(new_n1189), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1229), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1200), .B(new_n1228), .C1(new_n1164), .C2(new_n1189), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1255), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1271), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI211_X1 g1077(.A(KEYINPUT127), .B(new_n1255), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(G402));
endmodule


