//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G197gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT11), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  AND2_X1   g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G43gat), .A2(G50gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT15), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT14), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT14), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT89), .B(G36gat), .Z(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT90), .B(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT91), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n222), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n217), .B1(new_n227), .B2(new_n210), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT17), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  AOI211_X1 g028(.A(KEYINPUT15), .B(new_n208), .C1(new_n219), .C2(new_n220), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n210), .B1(new_n230), .B2(KEYINPUT91), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n218), .ZN(new_n232));
  INV_X1    g031(.A(new_n223), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n210), .B1(new_n233), .B2(new_n217), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G15gat), .B(G22gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G1gat), .ZN(new_n238));
  OAI21_X1  g037(.A(G8gat), .B1(new_n238), .B2(KEYINPUT92), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT16), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n237), .B1(new_n241), .B2(G1gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n236), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n232), .B(new_n234), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT93), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(KEYINPUT93), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n234), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(KEYINPUT94), .A3(new_n249), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n248), .B(KEYINPUT13), .Z(new_n260));
  INV_X1    g059(.A(KEYINPUT94), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT95), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n247), .A2(new_n249), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT18), .A3(new_n248), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n259), .A2(KEYINPUT95), .A3(new_n260), .A4(new_n262), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n202), .B(new_n207), .C1(new_n256), .C2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n207), .ZN(new_n271));
  INV_X1    g070(.A(new_n256), .ZN(new_n272));
  INV_X1    g071(.A(new_n269), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n207), .B1(new_n250), .B2(new_n251), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n265), .A2(new_n267), .A3(new_n275), .A4(new_n268), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT96), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n270), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G134gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G127gat), .B(G134gat), .Z(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(KEYINPUT1), .B2(new_n279), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT26), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n289), .A2(KEYINPUT26), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT27), .B(G183gat), .Z(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n297), .A2(new_n298), .A3(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT27), .B1(new_n291), .B2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(G183gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n303), .A3(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n300), .A2(new_n303), .A3(KEYINPUT70), .A4(new_n292), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n298), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n299), .B1(new_n308), .B2(KEYINPUT71), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n306), .A2(new_n310), .A3(new_n298), .A4(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n291), .A2(new_n292), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(new_n291), .B2(new_n292), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n322), .B2(KEYINPUT66), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT68), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n315), .A2(new_n316), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n318), .A2(new_n317), .B1(new_n291), .B2(new_n292), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(KEYINPUT66), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n287), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n331), .A2(KEYINPUT65), .A3(new_n333), .A4(new_n287), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n313), .A3(new_n320), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n330), .A2(new_n336), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n286), .B1(new_n312), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n291), .A2(KEYINPUT27), .ZN(new_n344));
  AOI21_X1  g143(.A(G190gat), .B1(new_n344), .B2(new_n301), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT70), .B1(new_n345), .B2(new_n300), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n307), .A2(new_n298), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT71), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n299), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n311), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n295), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n335), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n283), .A2(new_n285), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G227gat), .A2(G233gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(KEYINPUT64), .Z(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT34), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n356), .A3(KEYINPUT73), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n356), .A3(new_n357), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT34), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT34), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n312), .A2(new_n342), .A3(new_n286), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n355), .B1(new_n351), .B2(new_n354), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n358), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n358), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n343), .B2(new_n356), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n379), .B1(new_n382), .B2(KEYINPUT33), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n370), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n362), .A2(new_n363), .B1(new_n366), .B2(KEYINPUT72), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n385), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n369), .A4(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n391), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT36), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(KEYINPUT74), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G141gat), .B(G148gat), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT78), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  INV_X1    g207(.A(G148gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(G141gat), .ZN(new_n410));
  INV_X1    g209(.A(G141gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(G141gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n400), .A2(new_n405), .ZN(new_n415));
  NAND2_X1  g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n286), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n407), .A2(new_n418), .A3(KEYINPUT80), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT80), .B1(new_n407), .B2(new_n418), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n423), .B2(new_n286), .ZN(new_n424));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n398), .B(KEYINPUT5), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n418), .A3(KEYINPUT80), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n286), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n407), .A2(new_n418), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n355), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n425), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT4), .B1(new_n286), .B2(new_n419), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n355), .B1(new_n438), .B2(new_n431), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n428), .A2(KEYINPUT3), .A3(new_n429), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n355), .A2(new_n431), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n436), .A3(KEYINPUT81), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n437), .A2(new_n441), .A3(new_n425), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n435), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT5), .B1(new_n443), .B2(new_n436), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n441), .A3(new_n425), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT0), .ZN(new_n451));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  INV_X1    g254(.A(new_n453), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n456), .A3(new_n448), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n454), .A2(new_n460), .A3(new_n455), .A4(new_n457), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n446), .B2(new_n448), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G8gat), .B(G36gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(G226gat), .ZN(new_n468));
  INV_X1    g267(.A(G233gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT29), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n312), .B2(new_n342), .ZN(new_n473));
  XOR2_X1   g272(.A(G211gat), .B(G218gat), .Z(new_n474));
  XOR2_X1   g273(.A(G197gat), .B(G204gat), .Z(new_n475));
  AOI21_X1  g274(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT75), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(G197gat), .A2(G204gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(G197gat), .A2(G204gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n474), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n475), .A2(KEYINPUT75), .A3(new_n476), .ZN(new_n484));
  INV_X1    g283(.A(new_n474), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n470), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n351), .A2(new_n354), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n473), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT76), .B1(new_n483), .B2(new_n486), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n480), .A2(new_n481), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n485), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n482), .A2(new_n474), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n473), .B2(new_n489), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT30), .B(new_n467), .C1(new_n490), .C2(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n312), .A2(new_n342), .A3(new_n470), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n471), .B1(new_n351), .B2(new_n354), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n467), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n473), .A2(new_n489), .A3(new_n487), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n505), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT30), .B1(new_n510), .B2(new_n467), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n500), .A2(KEYINPUT77), .A3(new_n506), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n464), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n483), .B2(new_n486), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n431), .B1(new_n521), .B2(new_n438), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n487), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G228gat), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n522), .A2(new_n524), .B1(new_n525), .B2(new_n469), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n520), .C1(new_n419), .C2(KEYINPUT3), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n527), .A2(new_n491), .A3(new_n496), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT29), .B1(new_n493), .B2(new_n495), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n423), .B1(new_n531), .B2(KEYINPUT3), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(new_n469), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(G22gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n526), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n519), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G78gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n518), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n394), .A2(new_n397), .B1(new_n515), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n507), .A2(new_n511), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n439), .A2(new_n440), .B1(new_n443), .B2(new_n436), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(new_n425), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n453), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n424), .B2(new_n425), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n425), .B2(new_n551), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n554), .A2(KEYINPUT40), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT40), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n557), .A2(new_n558), .A3(new_n462), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n547), .B1(new_n550), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n510), .A2(new_n467), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n490), .B2(new_n499), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n473), .A2(new_n489), .A3(new_n498), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n501), .A2(new_n502), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT37), .B(new_n565), .C1(new_n566), .C2(new_n487), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .A4(new_n504), .ZN(new_n569));
  AND4_X1   g368(.A1(new_n458), .A2(new_n463), .A3(new_n562), .A4(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n503), .A2(KEYINPUT37), .A3(new_n505), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n504), .ZN(new_n573));
  INV_X1    g372(.A(new_n564), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n571), .A3(new_n504), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n570), .B1(new_n577), .B2(KEYINPUT87), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n579), .A2(new_n573), .A3(new_n574), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT87), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n580), .A2(new_n581), .A3(new_n568), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n560), .B(new_n561), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n580), .B2(new_n568), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n575), .A2(new_n576), .ZN(new_n586));
  INV_X1    g385(.A(new_n568), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT87), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n588), .A3(new_n570), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n561), .B1(new_n589), .B2(new_n560), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n548), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n458), .A2(KEYINPUT83), .B1(KEYINPUT6), .B2(new_n462), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n461), .B2(new_n594), .ZN(new_n595));
  AND4_X1   g394(.A1(new_n546), .A2(new_n387), .A3(new_n542), .A4(new_n391), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n387), .A2(new_n542), .A3(new_n546), .A4(new_n391), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n458), .A2(new_n463), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n592), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n598), .A2(new_n600), .A3(new_n550), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n278), .B1(new_n591), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  INV_X1    g404(.A(G71gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n537), .ZN(new_n607));
  XNOR2_X1  g406(.A(G57gat), .B(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT9), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n605), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G57gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(G64gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G57gat), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT98), .B1(new_n616), .B2(G64gat), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n611), .B2(G64gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n610), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT99), .Z(new_n622));
  XOR2_X1   g421(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n246), .B1(new_n620), .B2(new_n619), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n629), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n633), .A3(new_n627), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT7), .ZN(new_n641));
  NOR2_X1   g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(KEYINPUT8), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n229), .A2(new_n236), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n224), .A2(new_n228), .ZN(new_n650));
  INV_X1    g449(.A(new_n646), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n645), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n639), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n653), .A3(new_n639), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n656), .B1(new_n660), .B2(new_n654), .ZN(new_n661));
  XOR2_X1   g460(.A(G134gat), .B(G162gat), .Z(new_n662));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n659), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n664), .B(KEYINPUT101), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n659), .B2(new_n661), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n638), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n615), .A2(new_n618), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n645), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n647), .A2(new_n674), .A3(new_n610), .A4(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT102), .B1(new_n641), .B2(new_n644), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n652), .B1(new_n619), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT10), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n647), .A2(new_n619), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n673), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n677), .A2(new_n679), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(new_n673), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n683), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n687), .B(KEYINPUT104), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n673), .B(KEYINPUT105), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n681), .ZN(new_n695));
  INV_X1    g494(.A(new_n682), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n691), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n604), .A2(new_n672), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n464), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n550), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G8gat), .B1(new_n704), .B2(new_n549), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  MUX2_X1   g511(.A(new_n710), .B(new_n712), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g512(.A1(new_n394), .A2(new_n397), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n395), .A2(G15gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n704), .B2(new_n716), .ZN(G1326gat));
  INV_X1    g516(.A(new_n547), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT43), .B(G22gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  INV_X1    g520(.A(new_n278), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n659), .A2(new_n661), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n668), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n659), .A2(new_n661), .A3(new_n666), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n637), .A2(new_n726), .A3(new_n702), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n714), .B1(new_n718), .B2(new_n595), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n560), .B1(new_n578), .B2(new_n582), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(new_n583), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n722), .B(new_n727), .C1(new_n731), .C2(new_n602), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(G29gat), .A3(new_n464), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT45), .Z(new_n734));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n597), .B2(new_n601), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT35), .B1(new_n515), .B2(new_n598), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n596), .A2(new_n592), .A3(new_n599), .A4(new_n549), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n671), .B1(new_n731), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g542(.A(KEYINPUT44), .B(new_n671), .C1(new_n731), .C2(new_n602), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n637), .B(KEYINPUT107), .Z(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n278), .A3(new_n702), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n747), .B2(new_n464), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G29gat), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n747), .A2(KEYINPUT109), .A3(new_n464), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n734), .B1(new_n749), .B2(new_n750), .ZN(G1328gat));
  INV_X1    g550(.A(new_n215), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n732), .A2(new_n549), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT46), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n747), .B2(new_n549), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1329gat));
  NOR2_X1   g555(.A1(new_n395), .A2(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT47), .B1(new_n732), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n714), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n760), .A3(new_n744), .A4(new_n746), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n761), .B2(G43gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n764), .B(new_n759), .C1(new_n761), .C2(G43gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(G43gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(KEYINPUT110), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n732), .B2(new_n758), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n761), .B2(G43gat), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n763), .A2(new_n765), .B1(new_n768), .B2(new_n770), .ZN(G1330gat));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n547), .B1(new_n732), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT112), .B1(new_n604), .B2(new_n727), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n219), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n718), .A2(new_n219), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n747), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n775), .B(new_n779), .C1(new_n747), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1331gat));
  NAND3_X1  g580(.A1(new_n672), .A2(new_n278), .A3(new_n702), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n597), .A2(KEYINPUT108), .A3(new_n601), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n738), .B1(new_n736), .B2(new_n737), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n785), .B2(new_n591), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n706), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(new_n611), .Z(G1332gat));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n550), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT49), .B(G64gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1333gat));
  AOI21_X1  g591(.A(new_n606), .B1(new_n786), .B2(new_n760), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n395), .A2(G71gat), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n786), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n547), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g597(.A1(new_n722), .A2(new_n637), .A3(new_n703), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n726), .B1(new_n785), .B2(new_n591), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n744), .B(new_n799), .C1(new_n800), .C2(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n464), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n722), .A2(new_n637), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n671), .B(new_n803), .C1(new_n731), .C2(new_n740), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n591), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n671), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n464), .A2(new_n703), .A3(G85gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n802), .B1(new_n810), .B2(new_n811), .ZN(G1336gat));
  OAI21_X1  g611(.A(G92gat), .B1(new_n801), .B2(new_n549), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n703), .A2(G92gat), .A3(new_n549), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n818), .A3(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n813), .B(new_n817), .C1(new_n814), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT114), .B(G99gat), .Z(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n801), .B2(new_n714), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n703), .A2(new_n395), .A3(new_n823), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n810), .B2(new_n825), .ZN(G1338gat));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n718), .A2(new_n703), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT51), .B1(new_n800), .B2(new_n803), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n804), .A2(new_n805), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n517), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n718), .A2(new_n517), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n743), .A2(new_n744), .A3(new_n799), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n827), .A2(new_n828), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n830), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(G106gat), .B1(new_n809), .B2(new_n831), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n838), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(new_n829), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n840), .A2(new_n843), .ZN(G1339gat));
  NAND3_X1  g643(.A1(new_n672), .A2(new_n278), .A3(new_n703), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  INV_X1    g645(.A(new_n694), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n846), .B(new_n847), .C1(new_n680), .C2(new_n682), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n687), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n695), .A2(new_n696), .A3(new_n694), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n683), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n691), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n691), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT55), .B1(new_n849), .B2(new_n851), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n671), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n266), .A2(new_n248), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n260), .B1(new_n259), .B2(new_n262), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n206), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n276), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n863), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n702), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n278), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n864), .B1(new_n868), .B2(new_n726), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n845), .B1(new_n869), .B2(new_n745), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n598), .A2(new_n550), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n870), .A2(new_n706), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n722), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n870), .A2(new_n706), .A3(new_n549), .A4(new_n596), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT117), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n722), .A2(G113gat), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n875), .B2(new_n877), .ZN(G1340gat));
  AOI21_X1  g677(.A(G120gat), .B1(new_n872), .B2(new_n702), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n702), .A2(G120gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n875), .B2(new_n880), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n872), .A2(new_n882), .A3(new_n637), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n875), .A2(new_n745), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n882), .ZN(G1342gat));
  INV_X1    g684(.A(G134gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n872), .A2(new_n886), .A3(new_n671), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n875), .A2(new_n671), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n886), .ZN(G1343gat));
  NOR3_X1   g690(.A1(new_n760), .A2(new_n464), .A3(new_n550), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n870), .B2(new_n547), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n853), .A2(new_n857), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n270), .C1(new_n274), .C2(new_n277), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n671), .B1(new_n896), .B2(new_n866), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n638), .B1(new_n897), .B2(new_n864), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n894), .B(new_n718), .C1(new_n898), .C2(new_n845), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n892), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G141gat), .B1(new_n900), .B2(new_n278), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n870), .A2(new_n706), .A3(new_n547), .A4(new_n714), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n549), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n722), .A2(new_n411), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n901), .B(new_n902), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n903), .A2(new_n550), .A3(new_n907), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n892), .C1(new_n893), .C2(new_n899), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n722), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n913), .B2(G141gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n908), .B1(new_n914), .B2(new_n902), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n856), .A2(new_n858), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT116), .B1(new_n852), .B2(new_n691), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(new_n726), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n863), .B1(new_n918), .B2(KEYINPUT120), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n859), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n897), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n845), .B1(new_n922), .B2(new_n637), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n718), .B1(new_n923), .B2(KEYINPUT121), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n925), .B(new_n845), .C1(new_n922), .C2(new_n637), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n718), .A2(new_n894), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n870), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n702), .B(new_n892), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n904), .A2(new_n549), .A3(new_n905), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n703), .A2(G148gat), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n910), .A2(new_n912), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n409), .B1(new_n936), .B2(new_n702), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n937), .B2(KEYINPUT59), .ZN(G1345gat));
  NAND3_X1  g737(.A1(new_n910), .A2(new_n745), .A3(new_n912), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G155gat), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n638), .A2(G155gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n906), .B2(new_n941), .ZN(G1346gat));
  AOI21_X1  g741(.A(G162gat), .B1(new_n933), .B2(new_n671), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n671), .A2(G162gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n936), .B2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n706), .A2(new_n549), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n870), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n596), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n722), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(G169gat), .ZN(G1348gat));
  NAND4_X1  g749(.A1(new_n947), .A2(new_n718), .A3(new_n392), .A4(new_n702), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(G176gat), .ZN(G1349gat));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n638), .A2(new_n297), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n870), .A2(new_n596), .A3(new_n946), .A4(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n947), .A2(new_n596), .A3(new_n745), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G183gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n953), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n953), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT124), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n960), .A2(new_n963), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(G1350gat));
  XNOR2_X1  g766(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n948), .A2(new_n671), .B1(new_n292), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n292), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT126), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n969), .B(new_n971), .ZN(G1351gat));
  NAND2_X1  g771(.A1(new_n714), .A2(new_n946), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n870), .A2(new_n547), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n722), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n924), .A2(new_n926), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n894), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n973), .B1(new_n978), .B2(new_n929), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n722), .A2(G197gat), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(G1352gat));
  INV_X1    g781(.A(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n975), .A2(new_n983), .A3(new_n702), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  AND2_X1   g784(.A1(new_n979), .A2(new_n702), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n983), .ZN(G1353gat));
  INV_X1    g786(.A(G211gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n975), .A2(new_n988), .A3(new_n637), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n637), .B(new_n974), .C1(new_n927), .C2(new_n930), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n988), .B1(KEYINPUT127), .B2(new_n991), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n990), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  INV_X1    g795(.A(G218gat), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n975), .A2(new_n997), .A3(new_n671), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n979), .A2(new_n671), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n997), .ZN(G1355gat));
endmodule


