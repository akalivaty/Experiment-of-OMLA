//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G190gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT68), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n209));
  AND4_X1   g008(.A1(KEYINPUT68), .A2(new_n204), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n202), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n207), .A2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT26), .B2(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(G226gat), .A2(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n232), .B2(new_n219), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n226), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n233), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n236), .A2(new_n237), .B1(new_n226), .B2(new_n239), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT25), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n234), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(KEYINPUT25), .B(new_n230), .C1(new_n232), .C2(new_n219), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n231), .A2(G169gat), .A3(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n220), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT25), .A4(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n228), .B(new_n229), .C1(new_n246), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n250), .A2(new_n255), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  INV_X1    g058(.A(new_n245), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n253), .B1(new_n244), .B2(KEYINPUT65), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n258), .A2(new_n262), .B1(new_n218), .B2(new_n227), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n229), .A2(KEYINPUT29), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n257), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n267));
  NAND2_X1  g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G204gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G197gat), .ZN(new_n272));
  INV_X1    g071(.A(G197gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G204gat), .ZN(new_n274));
  AND4_X1   g073(.A1(new_n267), .A2(new_n270), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G197gat), .B(G204gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n276), .B2(new_n270), .ZN(new_n277));
  XOR2_X1   g076(.A(G211gat), .B(G218gat), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n275), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n274), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n276), .A2(new_n267), .A3(new_n270), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT73), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n279), .B1(new_n275), .B2(new_n277), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n278), .A3(new_n284), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n290), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n257), .B(new_n295), .C1(new_n263), .C2(new_n265), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(KEYINPUT37), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n292), .A2(KEYINPUT87), .A3(KEYINPUT37), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT37), .B1(new_n292), .B2(new_n296), .ZN(new_n302));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT74), .ZN(new_n304));
  XOR2_X1   g103(.A(G64gat), .B(G92gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n302), .A2(KEYINPUT38), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n306), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n292), .B2(new_n296), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT37), .ZN(new_n311));
  INV_X1    g110(.A(new_n296), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n228), .B1(new_n246), .B2(new_n256), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n264), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n295), .B1(new_n314), .B2(new_n257), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n309), .A3(new_n297), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n317), .B2(KEYINPUT38), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G134gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G127gat), .ZN(new_n321));
  INV_X1    g120(.A(G127gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(G113gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(KEYINPUT69), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(G120gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n325), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(new_n324), .B1(new_n321), .B2(new_n323), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT70), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n324), .B1(new_n331), .B2(new_n328), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n323), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT69), .B1(new_n330), .B2(G120gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n331), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n341), .B(new_n342), .C1(new_n346), .C2(new_n325), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  INV_X1    g150(.A(G148gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n357));
  INV_X1    g156(.A(G155gat), .ZN(new_n358));
  INV_X1    g157(.A(G162gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  AND2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT76), .B(new_n364), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n355), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n353), .A2(new_n354), .ZN(new_n367));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT77), .A4(new_n350), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n364), .A2(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n355), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n348), .A2(new_n375), .A3(KEYINPUT80), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n338), .A2(new_n347), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n366), .A2(new_n374), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT4), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n334), .A2(new_n337), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n382), .A3(new_n374), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(KEYINPUT4), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n377), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n387), .A3(new_n374), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT5), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n385), .A2(KEYINPUT81), .A3(new_n390), .A4(new_n393), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n379), .A2(new_n398), .A3(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n379), .B2(new_n389), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n383), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n392), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n376), .B1(new_n348), .B2(new_n375), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n383), .A2(KEYINPUT4), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n390), .B(new_n391), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT5), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n397), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G1gat), .B(G29gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(KEYINPUT85), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  INV_X1    g216(.A(new_n412), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n406), .A3(new_n418), .A4(new_n397), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n412), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n319), .A2(new_n413), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(new_n390), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n392), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(KEYINPUT86), .A3(new_n392), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n401), .A2(new_n392), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT86), .B1(new_n425), .B2(new_n392), .ZN(new_n434));
  AOI211_X1 g233(.A(new_n427), .B(new_n391), .C1(new_n385), .C2(new_n390), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n414), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n310), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n312), .A2(new_n315), .A3(new_n306), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n310), .A2(KEYINPUT30), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT40), .A4(new_n414), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n439), .A2(new_n445), .A3(new_n416), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n388), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n291), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n287), .A2(new_n448), .A3(new_n289), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n287), .A2(KEYINPUT82), .A3(new_n448), .A4(new_n289), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n450), .B1(new_n455), .B2(new_n375), .ZN(new_n456));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n387), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n459), .B2(new_n379), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  AOI221_X4 g267(.A(G22gat), .B1(new_n450), .B2(new_n460), .C1(new_n456), .C2(new_n457), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n458), .B2(new_n461), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT31), .B(G50gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT83), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n467), .B2(new_n471), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n424), .A2(new_n447), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  INV_X1    g277(.A(new_n473), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n469), .A2(new_n470), .A3(new_n468), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n466), .B1(new_n463), .B2(new_n465), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n407), .A2(new_n412), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n419), .A2(new_n417), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n421), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n445), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n478), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n263), .A2(new_n378), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n313), .A2(new_n348), .ZN(new_n493));
  INV_X1    g292(.A(G227gat), .ZN(new_n494));
  INV_X1    g293(.A(G233gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n497), .B(KEYINPUT32), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n493), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n509));
  INV_X1    g308(.A(new_n496), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n507), .B1(new_n514), .B2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g314(.A(new_n513), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n504), .A3(new_n518), .A4(new_n506), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n507), .A2(new_n514), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n504), .A3(new_n506), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(KEYINPUT36), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n477), .A2(new_n491), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n482), .A2(new_n484), .A3(new_n520), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT35), .B1(new_n527), .B2(new_n490), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n420), .A2(new_n423), .A3(new_n413), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n443), .A2(new_n530), .A3(new_n444), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n523), .B2(new_n522), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n476), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G43gat), .B(G50gat), .Z(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  NOR3_X1   g339(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND4_X1   g343(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(KEYINPUT89), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(KEYINPUT89), .B2(new_n543), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n538), .B1(new_n547), .B2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(G85gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(KEYINPUT8), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  NAND4_X1  g358(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n562), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n550), .A2(new_n570), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT96), .ZN(new_n576));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577));
  NOR2_X1   g376(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n576), .B(new_n579), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT16), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(G1gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n584), .B(new_n585), .C1(G1gat), .C2(new_n582), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G8gat), .ZN(new_n587));
  XOR2_X1   g386(.A(G57gat), .B(G64gat), .Z(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n588), .A2(KEYINPUT95), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(KEYINPUT95), .B2(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(G71gat), .ZN(new_n593));
  INV_X1    g392(.A(G78gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT94), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  MUX2_X1   g394(.A(KEYINPUT94), .B(new_n595), .S(new_n590), .Z(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT9), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n590), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n592), .A2(new_n596), .B1(new_n588), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n587), .B1(new_n599), .B2(KEYINPUT21), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n600), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  INV_X1    g411(.A(new_n600), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n611), .B2(new_n614), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n581), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT99), .B(new_n581), .C1(new_n617), .C2(new_n619), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n552), .A3(new_n553), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n550), .A2(new_n587), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT18), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT93), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(KEYINPUT93), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n587), .B(new_n549), .Z(new_n635));
  XOR2_X1   g434(.A(new_n629), .B(KEYINPUT13), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT11), .ZN(new_n640));
  INV_X1    g439(.A(G169gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G197gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n632), .A2(new_n634), .A3(new_n637), .A4(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n570), .A2(new_n599), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n599), .A2(new_n563), .A3(new_n567), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n570), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n651), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  AND4_X1   g468(.A1(new_n535), .A2(new_n622), .A3(new_n623), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n488), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  INV_X1    g472(.A(new_n670), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n489), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT101), .ZN(new_n678));
  OAI21_X1  g477(.A(G8gat), .B1(new_n674), .B2(new_n489), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n678), .B(new_n680), .C1(KEYINPUT42), .C2(new_n681), .ZN(G1325gat));
  INV_X1    g481(.A(new_n524), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n674), .A2(G15gat), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n525), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(G15gat), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT102), .Z(G1326gat));
  NAND2_X1  g487(.A1(new_n478), .A2(new_n485), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(G1327gat));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n528), .A2(new_n696), .A3(new_n533), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n526), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n528), .B2(new_n533), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n695), .B(new_n580), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n534), .A2(KEYINPUT104), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n526), .A3(new_n697), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n695), .A4(new_n580), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n581), .B1(new_n526), .B2(new_n534), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(new_n695), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n617), .A2(new_n619), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(new_n669), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n488), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n706), .A2(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(G29gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n671), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(G1328gat));
  OAI21_X1  g516(.A(G36gat), .B1(new_n711), .B2(new_n489), .ZN(new_n718));
  INV_X1    g517(.A(G36gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(new_n719), .A3(new_n445), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT106), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1329gat));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n685), .A3(new_n710), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G43gat), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n713), .A2(new_n727), .A3(new_n524), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT107), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT107), .B(new_n731), .C1(new_n726), .C2(new_n728), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(G1330gat));
  OAI21_X1  g532(.A(G50gat), .B1(new_n711), .B2(new_n476), .ZN(new_n734));
  INV_X1    g533(.A(G50gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n713), .A2(new_n735), .A3(new_n690), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(KEYINPUT48), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n736), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n708), .A2(new_n690), .A3(new_n710), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g540(.A1(new_n622), .A2(new_n623), .A3(new_n649), .A4(new_n668), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n703), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n671), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT108), .B(G57gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1332gat));
  AOI21_X1  g546(.A(new_n489), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n749), .B(new_n750), .Z(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743), .B2(new_n525), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n683), .A2(G71gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n690), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  INV_X1    g557(.A(new_n709), .ZN(new_n759));
  INV_X1    g558(.A(new_n668), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n648), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n708), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n708), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n488), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n759), .A2(new_n648), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n703), .A2(new_n580), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n580), .A4(new_n768), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n671), .A2(new_n555), .A3(new_n668), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n767), .B1(new_n773), .B2(new_n774), .ZN(G1336gat));
  OAI21_X1  g574(.A(KEYINPUT112), .B1(new_n762), .B2(new_n489), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n708), .A2(new_n777), .A3(new_n445), .A4(new_n761), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(G92gat), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n668), .A2(new_n556), .A3(new_n445), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT110), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n771), .A2(new_n772), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n782), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n445), .A3(new_n765), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n766), .B2(new_n525), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n760), .A2(G99gat), .A3(new_n683), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT113), .Z(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n773), .B2(new_n796), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n762), .B2(new_n476), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n476), .A2(new_n760), .A3(G106gat), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n785), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n799), .B(KEYINPUT114), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n773), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n763), .A2(new_n690), .A3(new_n765), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(G1339gat));
  NAND2_X1  g606(.A1(new_n671), .A2(new_n489), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n622), .A2(new_n623), .A3(new_n649), .A4(new_n760), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n655), .A2(new_n656), .A3(new_n651), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n664), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n657), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n811), .A2(new_n814), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n665), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n811), .A2(new_n814), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n648), .B(new_n819), .C1(KEYINPUT55), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n628), .A2(new_n629), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n635), .A2(new_n636), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n643), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n668), .A2(new_n647), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n580), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n580), .A2(new_n647), .A3(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(KEYINPUT55), .B2(new_n820), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n709), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n808), .B1(new_n809), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n476), .A3(new_n520), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n330), .A3(new_n648), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n690), .A2(new_n683), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n837), .A2(new_n648), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n839), .B2(new_n330), .ZN(G1340gat));
  NAND2_X1  g639(.A1(new_n668), .A2(new_n326), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n837), .A2(new_n668), .A3(new_n838), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n326), .ZN(G1341gat));
  AND3_X1   g644(.A1(new_n837), .A2(new_n759), .A3(new_n838), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n759), .A2(new_n322), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n846), .A2(new_n322), .B1(new_n832), .B2(new_n847), .ZN(G1342gat));
  NOR3_X1   g647(.A1(new_n581), .A2(new_n527), .A3(G134gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n852), .A2(new_n853), .B1(KEYINPUT56), .B2(new_n850), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n837), .A2(new_n580), .A3(new_n838), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n320), .B2(new_n855), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n685), .A2(new_n808), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n825), .B(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n811), .A2(new_n863), .A3(new_n814), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n811), .B2(new_n814), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n819), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n648), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n819), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n860), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n829), .B1(new_n870), .B2(new_n581), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n809), .B1(new_n871), .B2(new_n759), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n690), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n809), .A2(new_n830), .ZN(new_n874));
  INV_X1    g673(.A(new_n476), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n858), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(G141gat), .A3(new_n648), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n876), .A2(new_n858), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n648), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n351), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n880), .A2(KEYINPUT58), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1344gat));
  NAND3_X1  g687(.A1(new_n881), .A2(new_n352), .A3(new_n668), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n352), .C1(new_n879), .C2(new_n668), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n857), .B(KEYINPUT124), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n872), .B2(new_n690), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n877), .B(new_n476), .C1(new_n809), .C2(new_n830), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n668), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n890), .B2(new_n896), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n358), .A3(new_n759), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n879), .A2(new_n759), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n358), .ZN(G1346gat));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n359), .A3(new_n580), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n879), .A2(new_n580), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n359), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n671), .A2(new_n489), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n874), .A2(new_n835), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n649), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT126), .Z(new_n907));
  NOR2_X1   g706(.A1(new_n527), .A2(new_n489), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT125), .Z(new_n909));
  AOI211_X1 g708(.A(new_n671), .B(new_n909), .C1(new_n809), .C2(new_n830), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n641), .A3(new_n648), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n911), .ZN(G1348gat));
  OAI21_X1  g711(.A(G176gat), .B1(new_n905), .B2(new_n760), .ZN(new_n913));
  INV_X1    g712(.A(G176gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n914), .A3(new_n668), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1349gat));
  OAI21_X1  g715(.A(G183gat), .B1(new_n905), .B2(new_n709), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n202), .A3(new_n759), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n905), .B2(new_n581), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT61), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n215), .A3(new_n580), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n525), .A2(new_n904), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n876), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n648), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n893), .A2(new_n894), .ZN(new_n928));
  INV_X1    g727(.A(new_n925), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n649), .A2(new_n273), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  OAI211_X1 g731(.A(new_n668), .B(new_n929), .C1(new_n893), .C2(new_n894), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n760), .A2(G204gat), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n874), .A2(new_n875), .A3(new_n929), .A4(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  INV_X1    g741(.A(G211gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n943), .A3(new_n759), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n759), .B(new_n929), .C1(new_n893), .C2(new_n894), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  INV_X1    g747(.A(G218gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n926), .A2(new_n949), .A3(new_n580), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n580), .A3(new_n929), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n949), .ZN(G1355gat));
endmodule


