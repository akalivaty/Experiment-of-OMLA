//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G141gat), .B(G148gat), .Z(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n210), .C1(new_n214), .C2(KEYINPUT2), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n212), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT29), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n208), .A2(new_n219), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G228gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n223), .B(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n226), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n223), .B(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(G22gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n227), .A2(new_n231), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G78gat), .B(G106gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT31), .B(G50gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n232), .A3(new_n239), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT70), .B(G120gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT71), .B(G113gat), .ZN(new_n247));
  INV_X1    g046(.A(G120gat), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n245), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(G113gat), .B2(G120gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n253), .B1(G113gat), .B2(G120gat), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n254), .A2(new_n251), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n216), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT4), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n216), .A2(new_n217), .ZN(new_n259));
  INV_X1    g058(.A(new_n256), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n218), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT5), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n256), .B(new_n216), .Z(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G1gat), .B(G29gat), .ZN(new_n272));
  INV_X1    g071(.A(G85gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n270), .B1(new_n266), .B2(new_n268), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(new_n264), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n281), .A2(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT6), .B1(new_n271), .B2(new_n277), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT82), .A3(new_n281), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n293), .B(KEYINPUT66), .Z(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT65), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT68), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n300), .B2(new_n301), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n309), .B(KEYINPUT67), .Z(new_n310));
  OAI211_X1 g109(.A(new_n297), .B(new_n299), .C1(new_n307), .C2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n302), .A3(new_n306), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n299), .A2(new_n296), .A3(new_n293), .A4(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n295), .B(KEYINPUT26), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n317), .A2(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT28), .B1(new_n319), .B2(new_n301), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n292), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(KEYINPUT77), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n323), .B(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n316), .ZN(new_n329));
  INV_X1    g128(.A(new_n292), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n326), .A2(new_n208), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(KEYINPUT29), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n329), .A2(new_n333), .B1(new_n324), .B2(new_n330), .ZN(new_n334));
  INV_X1    g133(.A(new_n208), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G64gat), .B(G92gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT78), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND3_X1  g139(.A1(new_n332), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT79), .B1(new_n341), .B2(KEYINPUT80), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n341), .B2(KEYINPUT79), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n332), .A2(new_n336), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n342), .A2(new_n344), .B1(new_n345), .B2(new_n340), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n342), .A2(KEYINPUT30), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n244), .B1(new_n291), .B2(new_n349), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n279), .A2(KEYINPUT86), .A3(new_n264), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT86), .B1(new_n279), .B2(new_n264), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n276), .B(KEYINPUT85), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n286), .B1(new_n288), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT37), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n340), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n357), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT38), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n326), .A2(new_n335), .A3(new_n327), .A4(new_n331), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n334), .B2(new_n208), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT38), .B(new_n340), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n356), .A2(new_n362), .A3(new_n341), .A4(new_n366), .ZN(new_n367));
  OR3_X1    g166(.A1(new_n262), .A2(KEYINPUT39), .A3(new_n263), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n262), .A2(new_n263), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n267), .A2(new_n263), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT39), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n368), .B(new_n353), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT40), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n355), .B(new_n373), .C1(new_n346), .C2(new_n347), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n243), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G227gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n256), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n329), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n378), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT75), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n383), .B2(new_n386), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n378), .A3(new_n382), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n397), .B(KEYINPUT32), .C1(new_n398), .C2(new_n396), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n390), .A2(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n402), .A3(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(KEYINPUT36), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT76), .B1(new_n393), .B2(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n406), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT76), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(KEYINPUT36), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n350), .A2(new_n375), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n243), .A2(new_n404), .A3(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n243), .A2(new_n404), .A3(KEYINPUT87), .A4(new_n406), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n290), .A2(new_n415), .A3(new_n348), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT88), .B1(new_n417), .B2(KEYINPUT35), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(new_n243), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n356), .A2(KEYINPUT35), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n419), .A2(new_n420), .A3(new_n349), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n412), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G43gat), .B(G50gat), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n426));
  NAND2_X1  g225(.A1(G29gat), .A2(G36gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n427), .B(KEYINPUT91), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n429));
  OR3_X1    g228(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(KEYINPUT90), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n427), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(G1gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(G1gat), .B2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(G8gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n438), .A2(new_n439), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n438), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n452), .A3(new_n450), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n446), .B(new_n438), .Z(new_n457));
  XOR2_X1   g256(.A(new_n452), .B(KEYINPUT13), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n453), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G169gat), .B(G197gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT12), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n453), .A2(new_n466), .A3(new_n456), .A4(new_n459), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n424), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G57gat), .B(G64gat), .Z(new_n473));
  OR2_X1    g272(.A1(G71gat), .A2(G78gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(G71gat), .A2(G78gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G57gat), .B(G64gat), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n475), .B(new_n474), .C1(new_n480), .C2(new_n477), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT93), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT21), .ZN(new_n487));
  INV_X1    g286(.A(new_n482), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n488), .A2(KEYINPUT21), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n449), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n449), .B2(new_n489), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n492));
  XNOR2_X1  g291(.A(G183gat), .B(G211gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n491), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT92), .ZN(new_n497));
  XNOR2_X1  g296(.A(G127gat), .B(G155gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504));
  INV_X1    g303(.A(G92gat), .ZN(new_n505));
  AOI22_X1  g304(.A1(KEYINPUT8), .A2(new_n504), .B1(new_n273), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n504), .ZN(new_n511));
  NOR2_X1   g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G99gat), .ZN(new_n515));
  INV_X1    g314(.A(G106gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT95), .B1(new_n517), .B2(new_n504), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n506), .B(new_n510), .C1(new_n514), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT8), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n273), .A2(new_n505), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n507), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n513), .B1(new_n511), .B2(new_n512), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n517), .A2(KEYINPUT95), .A3(new_n504), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n503), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n525), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT96), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n438), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n440), .A2(new_n447), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(new_n533), .ZN(new_n537));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT94), .ZN(new_n541));
  XOR2_X1   g340(.A(G134gat), .B(G162gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n502), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT99), .ZN(new_n551));
  XNOR2_X1  g350(.A(G120gat), .B(G148gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n529), .A2(new_n488), .A3(new_n532), .ZN(new_n554));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n482), .B1(new_n519), .B2(new_n528), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n557), .B2(KEYINPUT98), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n532), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n482), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n556), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT10), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n484), .B2(new_n485), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n567), .A2(new_n533), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n555), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n557), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n558), .B1(new_n571), .B2(KEYINPUT98), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n553), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n549), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n472), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT100), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n291), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G1gat), .ZN(G1324gat));
  INV_X1    g379(.A(KEYINPUT42), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT101), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT16), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n349), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G8gat), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n578), .A2(new_n445), .A3(new_n349), .A4(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n349), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n581), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G1325gat));
  AOI21_X1  g388(.A(G15gat), .B1(new_n578), .B2(new_n410), .ZN(new_n590));
  INV_X1    g389(.A(new_n411), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(G15gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n578), .B2(new_n592), .ZN(G1326gat));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n244), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT43), .B(G22gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(G1327gat));
  INV_X1    g395(.A(new_n502), .ZN(new_n597));
  INV_X1    g396(.A(new_n548), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n574), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT102), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n472), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G29gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n291), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT45), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n574), .B(KEYINPUT103), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n606), .A2(new_n471), .A3(new_n502), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT44), .B1(new_n424), .B2(new_n548), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610));
  INV_X1    g409(.A(new_n423), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n611), .A2(new_n418), .A3(new_n421), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n610), .B(new_n598), .C1(new_n612), .C2(new_n412), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(new_n291), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n604), .B1(new_n615), .B2(new_n602), .ZN(G1328gat));
  NOR2_X1   g415(.A1(new_n348), .A2(G36gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n472), .A2(new_n600), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n609), .A2(new_n613), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n621), .A2(KEYINPUT105), .A3(new_n349), .A4(new_n607), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G36gat), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT105), .B1(new_n614), .B2(new_n349), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT106), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT106), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n620), .B(new_n627), .C1(new_n623), .C2(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(G1329gat));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n591), .ZN(new_n630));
  INV_X1    g429(.A(G43gat), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n410), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n630), .A2(G43gat), .B1(new_n601), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g433(.A(KEYINPUT107), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n614), .A2(new_n244), .ZN(new_n636));
  INV_X1    g435(.A(G50gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n601), .A2(new_n637), .A3(new_n244), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT48), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI221_X1 g441(.A(new_n639), .B1(new_n635), .B2(KEYINPUT48), .C1(new_n636), .C2(new_n637), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(G1331gat));
  NOR4_X1   g443(.A1(new_n424), .A2(new_n470), .A3(new_n549), .A4(new_n605), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n291), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g446(.A(new_n348), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT108), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1333gat));
  INV_X1    g451(.A(G71gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n645), .B2(new_n591), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n410), .A2(new_n653), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n645), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g456(.A1(new_n645), .A2(new_n244), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G78gat), .ZN(G1335gat));
  INV_X1    g458(.A(new_n621), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n502), .A2(new_n470), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n575), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT109), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n660), .A2(new_n290), .A3(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n598), .B(new_n661), .C1(new_n612), .C2(new_n412), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT51), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n422), .A2(new_n423), .ZN(new_n669));
  INV_X1    g468(.A(new_n412), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n598), .A4(new_n661), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n291), .A2(new_n273), .A3(new_n575), .ZN(new_n675));
  OAI22_X1  g474(.A1(new_n665), .A2(new_n273), .B1(new_n674), .B2(new_n675), .ZN(G1336gat));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n666), .A2(new_n677), .A3(new_n667), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n348), .A2(G92gat), .A3(new_n605), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n678), .B(new_n679), .C1(new_n673), .C2(new_n677), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n348), .B(new_n664), .C1(new_n609), .C2(new_n613), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n505), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT52), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT52), .B1(new_n673), .B2(new_n679), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n685));
  OAI21_X1  g484(.A(G92gat), .B1(new_n681), .B2(KEYINPUT111), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(G1337gat));
  NOR3_X1   g487(.A1(new_n660), .A2(new_n411), .A3(new_n664), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n410), .A2(new_n515), .A3(new_n575), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n689), .A2(new_n515), .B1(new_n674), .B2(new_n690), .ZN(G1338gat));
  NOR3_X1   g490(.A1(new_n243), .A2(G106gat), .A3(new_n605), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n678), .B(new_n692), .C1(new_n673), .C2(new_n677), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n621), .A2(new_n244), .A3(new_n663), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G106gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT53), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n673), .A2(new_n692), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1339gat));
  INV_X1    g500(.A(new_n555), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n566), .B1(new_n554), .B2(new_n556), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n567), .A2(new_n533), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n553), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n702), .A3(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n569), .A2(KEYINPUT54), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(KEYINPUT55), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT114), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n707), .A2(new_n709), .A3(new_n712), .A4(KEYINPUT55), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n572), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n707), .A2(new_n709), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT55), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND4_X1   g517(.A1(KEYINPUT115), .A2(new_n714), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n572), .B1(new_n711), .B2(new_n713), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT115), .B1(new_n720), .B2(new_n718), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n470), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n451), .A2(new_n452), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n457), .A2(new_n458), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n465), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n469), .A2(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n726), .A2(KEYINPUT116), .A3(new_n574), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT116), .B1(new_n726), .B2(new_n574), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n598), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n718), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n720), .A2(KEYINPUT115), .A3(new_n718), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n548), .A2(new_n726), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT117), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n727), .A2(new_n728), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n735), .B2(new_n470), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n739), .B(new_n740), .C1(new_n742), .C2(new_n598), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n743), .A3(new_n597), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n576), .A2(new_n471), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n744), .A2(KEYINPUT118), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT118), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n419), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n349), .A2(new_n290), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G113gat), .B1(new_n754), .B2(new_n471), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n748), .A2(new_n415), .A3(new_n416), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n751), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n471), .A2(new_n247), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(G1340gat));
  OAI21_X1  g558(.A(G120gat), .B1(new_n754), .B2(new_n605), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n574), .A2(new_n246), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT119), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n757), .B2(new_n762), .ZN(G1341gat));
  NAND3_X1  g562(.A1(new_n756), .A2(new_n502), .A3(new_n751), .ZN(new_n764));
  INV_X1    g563(.A(G127gat), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n597), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n764), .A2(new_n765), .B1(new_n753), .B2(new_n766), .ZN(G1342gat));
  OR3_X1    g566(.A1(new_n757), .A2(G134gat), .A3(new_n548), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(KEYINPUT56), .ZN(new_n769));
  OAI21_X1  g568(.A(G134gat), .B1(new_n754), .B2(new_n548), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(KEYINPUT56), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(G1343gat));
  NOR2_X1   g571(.A1(new_n726), .A2(new_n574), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT55), .B1(new_n716), .B2(KEYINPUT121), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT121), .B2(new_n716), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n720), .A3(new_n470), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n598), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT122), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n737), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(KEYINPUT122), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n502), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n745), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n244), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n591), .B(new_n752), .C1(new_n785), .C2(KEYINPUT57), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n746), .A2(new_n747), .A3(new_n243), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G141gat), .B1(new_n790), .B2(new_n471), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n411), .A3(new_n751), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n471), .A2(G141gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g594(.A(G148gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n752), .A2(new_n591), .A3(new_n574), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n787), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT123), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n748), .A2(new_n800), .A3(KEYINPUT57), .A4(new_n244), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n744), .A2(new_n745), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n744), .A2(KEYINPUT118), .A3(new_n745), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n804), .A2(KEYINPUT57), .A3(new_n244), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT123), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n731), .A2(new_n548), .A3(new_n726), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n597), .B1(new_n779), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n745), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n788), .B1(new_n810), .B2(new_n243), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n801), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n797), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n796), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT124), .A3(new_n797), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n799), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n790), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT59), .B(new_n796), .C1(new_n818), .C2(new_n575), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n798), .B1(new_n817), .B2(new_n819), .ZN(G1345gat));
  INV_X1    g619(.A(G155gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n790), .A2(new_n821), .A3(new_n597), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n792), .A2(new_n597), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(G1346gat));
  OAI21_X1  g623(.A(G162gat), .B1(new_n790), .B2(new_n548), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n548), .A2(G162gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n792), .B2(new_n826), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n291), .A2(new_n348), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n756), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G169gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n470), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n748), .A2(new_n749), .A3(new_n828), .ZN(new_n832));
  OAI21_X1  g631(.A(G169gat), .B1(new_n832), .B2(new_n471), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1348gat));
  INV_X1    g633(.A(G176gat), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n832), .A2(new_n835), .A3(new_n605), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n829), .A2(new_n575), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n835), .ZN(G1349gat));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n319), .A3(new_n502), .ZN(new_n839));
  OAI21_X1  g638(.A(G183gat), .B1(new_n832), .B2(new_n597), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g641(.A1(new_n832), .A2(new_n548), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n843), .A2(KEYINPUT125), .A3(new_n301), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT125), .B1(new_n843), .B2(new_n301), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n301), .A3(new_n598), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(KEYINPUT61), .A3(new_n845), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1351gat));
  AND2_X1   g650(.A1(new_n828), .A2(new_n411), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n812), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G197gat), .B1(new_n853), .B2(new_n471), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n787), .A2(new_n852), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n855), .A2(G197gat), .A3(new_n471), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1352gat));
  NOR3_X1   g656(.A1(new_n855), .A2(G204gat), .A3(new_n574), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT62), .ZN(new_n859));
  OAI21_X1  g658(.A(G204gat), .B1(new_n853), .B2(new_n605), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1353gat));
  NAND3_X1  g660(.A1(new_n812), .A2(new_n502), .A3(new_n852), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT63), .B1(new_n862), .B2(G211gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n502), .A2(new_n203), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n863), .A2(new_n864), .B1(new_n855), .B2(new_n865), .ZN(G1354gat));
  OAI21_X1  g665(.A(new_n204), .B1(new_n855), .B2(new_n548), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT126), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT126), .ZN(new_n869));
  INV_X1    g668(.A(new_n853), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n548), .A2(new_n204), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT127), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n872), .ZN(G1355gat));
endmodule


