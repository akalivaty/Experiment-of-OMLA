//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n210), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n202), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n215), .B1(KEYINPUT1), .B2(new_n224), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n210), .A2(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT74), .B(KEYINPUT11), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT75), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(KEYINPUT75), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n209), .A2(G20), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g0062(.A(new_n254), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n268));
  OR3_X1    g0068(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(G68), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n259), .A2(new_n260), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n225), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n281), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(new_n279), .A3(G232), .A4(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT73), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n275), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT68), .B1(new_n273), .B2(new_n225), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n293), .A2(new_n294), .A3(G1), .A4(G13), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G238), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT67), .A2(G45), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT67), .A2(G45), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n302), .A2(new_n292), .A3(new_n295), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n290), .A2(new_n291), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT13), .B1(new_n289), .B2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(G169), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n310), .B2(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n272), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(G200), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n308), .A2(G190), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n271), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n322), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT8), .A2(G58), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT70), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n326), .B1(new_n331), .B2(KEYINPUT8), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n210), .A3(G33), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n263), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n264), .ZN(new_n336));
  INV_X1    g0136(.A(G50), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n266), .B2(new_n337), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n335), .A2(KEYINPUT9), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT9), .B1(new_n335), .B2(new_n339), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n296), .A2(G226), .A3(new_n297), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G222), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G223), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n286), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n274), .C1(G77), .C2(new_n286), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n348), .A3(new_n305), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n342), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n324), .B(new_n325), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n281), .A2(G232), .B1(G107), .B2(new_n280), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n286), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n216), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n274), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n296), .A2(G244), .A3(new_n297), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(new_n305), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(G179), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n264), .A2(G77), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n266), .A2(new_n250), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT8), .B(G58), .Z(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n251), .B2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n364), .B(new_n365), .C1(new_n254), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(G169), .B1(new_n359), .B2(new_n361), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n363), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(G200), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n370), .C1(new_n374), .C2(new_n362), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n352), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n377), .A2(KEYINPUT72), .A3(KEYINPUT10), .A4(new_n353), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n335), .A2(new_n339), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n350), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G169), .B2(new_n350), .ZN(new_n382));
  AND4_X1   g0182(.A1(new_n355), .A2(new_n376), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n286), .B2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT78), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n280), .A2(new_n390), .A3(new_n210), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n217), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n248), .A2(G159), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n202), .B1(new_n331), .B2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n210), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n384), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT70), .B(G58), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n228), .B1(new_n398), .B2(new_n217), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n276), .A2(KEYINPUT77), .A3(G33), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n286), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n388), .B1(new_n403), .B2(new_n210), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n277), .A2(new_n279), .A3(new_n402), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n276), .A2(KEYINPUT77), .A3(G33), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n388), .A3(new_n210), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT16), .B(new_n400), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT79), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n384), .C1(new_n392), .C2(new_n395), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n397), .A2(new_n254), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n332), .A2(new_n336), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n266), .B2(new_n332), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT80), .ZN(new_n417));
  INV_X1    g0217(.A(G169), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n406), .ZN(new_n419));
  INV_X1    g0219(.A(G226), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G223), .B2(G1698), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G87), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n278), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n275), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n292), .A2(G232), .A3(new_n295), .A4(new_n297), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n305), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n418), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n305), .A2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n422), .B1(new_n406), .B2(new_n405), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n274), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n434), .A3(new_n380), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n417), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n417), .A3(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT18), .B1(new_n416), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n431), .A2(new_n417), .A3(new_n435), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n436), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n412), .A2(new_n415), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n428), .A2(G190), .A3(new_n430), .ZN(new_n446));
  AOI21_X1  g0246(.A(G200), .B1(new_n432), .B2(new_n434), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n351), .B1(new_n428), .B2(new_n430), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n432), .A2(new_n434), .A3(new_n374), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT81), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n412), .B(new_n415), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n448), .B1(new_n446), .B2(new_n447), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(KEYINPUT17), .A3(new_n415), .A4(new_n412), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n440), .A2(new_n445), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n316), .A2(new_n319), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND4_X1   g0264(.A1(new_n320), .A2(new_n383), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT86), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n296), .A2(G257), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n467), .A2(new_n303), .A3(G1), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n292), .A2(new_n473), .A3(new_n474), .A4(new_n295), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G244), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1698), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n286), .A2(KEYINPUT4), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n419), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n479), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n405), .B2(new_n406), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n483), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n274), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n476), .B1(new_n492), .B2(KEYINPUT85), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n494), .A3(new_n274), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n351), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n476), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(G190), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n206), .B1(new_n387), .B2(new_n391), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n248), .A2(G77), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT82), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n205), .B2(G107), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n207), .A2(new_n503), .A3(new_n505), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n500), .B(new_n501), .C1(new_n210), .C2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n254), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n336), .A2(new_n205), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n209), .A2(G33), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n263), .A2(new_n264), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n205), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n498), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n466), .B1(new_n496), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT4), .B1(new_n489), .B2(new_n484), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT84), .B1(new_n403), .B2(new_n488), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n482), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT85), .B1(new_n523), .B2(new_n275), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n495), .A2(new_n524), .A3(new_n497), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n501), .B1(new_n510), .B2(new_n210), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(KEYINPUT83), .B2(new_n499), .ZN(new_n528));
  INV_X1    g0328(.A(new_n512), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n263), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT86), .A4(new_n498), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n493), .A2(KEYINPUT87), .A3(new_n380), .A4(new_n495), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n495), .A2(new_n524), .A3(new_n380), .A4(new_n497), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n476), .B1(new_n491), .B2(new_n274), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n530), .A2(new_n517), .B1(new_n538), .B2(G169), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n520), .A2(new_n532), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(G238), .A2(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n478), .A2(G1698), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n405), .B2(new_n406), .ZN(new_n545));
  AND2_X1   g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n274), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G250), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n468), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n296), .B1(new_n474), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT88), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G190), .A3(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(G20), .B(new_n217), .C1(new_n405), .C2(new_n406), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n251), .B2(new_n205), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT89), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT89), .B(new_n557), .C1(new_n251), .C2(new_n205), .ZN(new_n561));
  NAND3_X1  g0361(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n210), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(G87), .B2(new_n207), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n254), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n368), .A2(new_n336), .ZN(new_n567));
  INV_X1    g0367(.A(new_n516), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G87), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT88), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT88), .B1(new_n547), .B2(new_n550), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n555), .B(new_n571), .C1(new_n574), .C2(new_n351), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n553), .A2(new_n380), .A3(new_n554), .ZN(new_n576));
  XOR2_X1   g0376(.A(new_n368), .B(KEYINPUT90), .Z(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n568), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n566), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n579), .C1(new_n574), .C2(G169), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(KEYINPUT22), .A2(G87), .ZN(new_n582));
  AOI211_X1 g0382(.A(G20), .B(new_n582), .C1(new_n405), .C2(new_n406), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n210), .A2(G87), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n280), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT23), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n210), .B2(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(new_n210), .B2(new_n546), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT24), .B1(new_n583), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n582), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n419), .A2(new_n210), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n586), .A4(new_n590), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n254), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n264), .A2(new_n599), .A3(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n264), .B2(G107), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n568), .A2(G107), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n548), .A2(new_n345), .ZN(new_n605));
  INV_X1    g0405(.A(G257), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G1698), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n405), .B2(new_n406), .ZN(new_n609));
  INV_X1    g0409(.A(G294), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n278), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n274), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n471), .A2(new_n292), .A3(G264), .A4(new_n295), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT92), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(KEYINPUT92), .A3(new_n613), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n475), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n351), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(new_n374), .A3(new_n475), .A4(new_n613), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT93), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n604), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n616), .A2(G179), .A3(new_n475), .A4(new_n617), .ZN(new_n623));
  INV_X1    g0423(.A(new_n475), .ZN(new_n624));
  OAI21_X1  g0424(.A(G169), .B1(new_n614), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(new_n625), .B1(new_n598), .B2(new_n603), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n345), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(G264), .B2(new_n345), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n406), .B2(new_n405), .ZN(new_n631));
  XNOR2_X1  g0431(.A(KEYINPUT91), .B(G303), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n286), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n274), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n471), .A2(new_n292), .A3(G270), .A4(new_n295), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n475), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n636), .A3(G190), .ZN(new_n637));
  INV_X1    g0437(.A(G116), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n253), .A2(new_n225), .B1(G20), .B2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n481), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(KEYINPUT20), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT20), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n336), .A2(new_n638), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n516), .B2(new_n638), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n635), .A2(new_n475), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n403), .A2(new_n630), .B1(new_n286), .B2(new_n632), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n274), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n637), .B(new_n646), .C1(new_n649), .C2(new_n351), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  OAI21_X1  g0451(.A(G169), .B1(new_n643), .B2(new_n645), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n634), .A2(new_n636), .ZN(new_n654));
  OAI221_X1 g0454(.A(new_n644), .B1(new_n516), .B2(new_n638), .C1(new_n641), .C2(new_n642), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT21), .A4(G169), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n655), .A3(G179), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n650), .A2(new_n653), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n628), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n465), .A2(new_n541), .A3(new_n581), .A4(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n382), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n440), .A2(new_n445), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n310), .A2(G169), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n313), .A3(new_n312), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n363), .A2(new_n370), .A3(new_n371), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n665), .A2(new_n272), .B1(new_n319), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n455), .A2(new_n459), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT95), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n378), .A2(new_n355), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n661), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n551), .A2(new_n418), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n576), .A2(new_n579), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT94), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n570), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n551), .A2(G200), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n555), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n626), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n683), .A3(new_n622), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n520), .A2(new_n532), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n537), .A2(new_n540), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n581), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT26), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n539), .B1(new_n533), .B2(new_n536), .ZN(new_n690));
  INV_X1    g0490(.A(new_n681), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n687), .A2(new_n676), .A3(new_n689), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n465), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n674), .A2(new_n695), .ZN(G369));
  NAND3_X1  g0496(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n700));
  INV_X1    g0500(.A(G213), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT97), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n704), .A2(G343), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n604), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT98), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n710), .A2(new_n627), .B1(new_n626), .B2(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n655), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n682), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n658), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n707), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n682), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n710), .A2(new_n627), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n626), .A2(new_n719), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n213), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n229), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n676), .B(KEYINPUT100), .Z(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n687), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT26), .B1(new_n686), .B2(new_n681), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n690), .A2(new_n692), .A3(new_n581), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n719), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n692), .B1(new_n690), .B2(new_n581), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n686), .A2(new_n681), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n692), .ZN(new_n741));
  INV_X1    g0541(.A(new_n676), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n541), .B2(new_n684), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n707), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n738), .B1(new_n744), .B2(KEYINPUT29), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n612), .A2(KEYINPUT92), .A3(new_n613), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT92), .B1(new_n612), .B2(new_n613), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n634), .A2(new_n636), .A3(G179), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n538), .A2(new_n574), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n572), .A2(new_n749), .A3(new_n573), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n748), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n654), .A2(new_n551), .A3(new_n380), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n748), .B2(new_n475), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n525), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT31), .B1(new_n759), .B2(new_n707), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT99), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n707), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT99), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n622), .A2(new_n626), .A3(new_n658), .A4(new_n707), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n685), .A2(new_n686), .A3(new_n581), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n762), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n745), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT101), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT101), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n745), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n731), .B1(new_n777), .B2(G1), .ZN(G364));
  AND2_X1   g0578(.A1(new_n210), .A2(G13), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n209), .B1(new_n779), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n726), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n725), .A2(new_n419), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n299), .A2(new_n301), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n784), .B1(new_n229), .B2(new_n785), .C1(new_n246), .C2(new_n467), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n213), .A2(new_n286), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(G116), .B2(new_n213), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT102), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n225), .B1(G20), .B2(new_n418), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(G20), .A2(G179), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT103), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n374), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n800), .A2(new_n250), .B1(new_n802), .B2(new_n337), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n798), .A2(new_n351), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G68), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n210), .A2(G179), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(new_n374), .A3(new_n351), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  OR3_X1    g0608(.A1(new_n807), .A2(KEYINPUT32), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G87), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n807), .B2(new_n808), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n374), .A3(G200), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G107), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n210), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n205), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n817), .A2(new_n280), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n797), .A2(G190), .A3(new_n351), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n822), .A2(KEYINPUT104), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(KEYINPUT104), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n805), .B(new_n821), .C1(new_n398), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n819), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n801), .A2(G326), .B1(G294), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n800), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT105), .Z(new_n831));
  INV_X1    g0631(.A(new_n807), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n286), .B1(new_n832), .B2(G329), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  INV_X1    g0634(.A(G303), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n814), .C1(new_n835), .C2(new_n810), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT106), .B(KEYINPUT33), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(G317), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n804), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G322), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n825), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n826), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n783), .B(new_n795), .C1(new_n842), .C2(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n792), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n715), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n782), .B1(new_n715), .B2(G330), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G330), .B2(new_n715), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  AOI211_X1 g0649(.A(new_n286), .B(new_n820), .C1(G311), .C2(new_n832), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n425), .B2(new_n814), .C1(new_n206), .C2(new_n810), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G303), .B2(new_n801), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G116), .A2(new_n799), .B1(new_n804), .B2(G283), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n610), .C2(new_n825), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n819), .A2(new_n398), .B1(new_n814), .B2(new_n217), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n419), .B1(new_n856), .B2(new_n807), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G50), .C2(new_n811), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n799), .A2(G159), .B1(new_n801), .B2(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  INV_X1    g0660(.A(new_n804), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT107), .B(G143), .Z(new_n862));
  OAI221_X1 g0662(.A(new_n859), .B1(new_n860), .B2(new_n861), .C1(new_n825), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT34), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n863), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(KEYINPUT34), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n854), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT108), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n793), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n375), .B1(new_n370), .B2(new_n719), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n372), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n666), .A2(new_n719), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(new_n791), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n793), .A2(new_n790), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n783), .B1(new_n250), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n870), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n376), .A2(new_n719), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n694), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT109), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n744), .A2(new_n884), .A3(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n694), .A2(new_n719), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT109), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(new_n772), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n782), .B1(new_n888), .B2(new_n772), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n880), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  AND2_X1   g0692(.A1(new_n704), .A2(new_n706), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n662), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n409), .A2(new_n254), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n400), .B1(new_n404), .B2(new_n408), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT16), .B1(new_n896), .B2(KEYINPUT111), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT111), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(new_n400), .C1(new_n404), .C2(new_n408), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n893), .B1(new_n900), .B2(new_n414), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n460), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n414), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n901), .B(new_n453), .C1(new_n904), .C2(new_n439), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n442), .A2(new_n443), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n443), .A2(new_n893), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n453), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n903), .B2(new_n911), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n271), .A2(new_n317), .A3(new_n318), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n272), .B(new_n707), .C1(new_n665), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n272), .A2(new_n707), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n316), .A2(new_n319), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n881), .B1(new_n741), .B2(new_n743), .ZN(new_n921));
  INV_X1    g0721(.A(new_n873), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n903), .A2(new_n911), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n907), .A2(new_n908), .A3(new_n453), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT112), .B1(new_n929), .B2(new_n910), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n908), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n460), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(KEYINPUT112), .A3(new_n910), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n913), .B1(new_n935), .B2(new_n925), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n927), .B1(new_n936), .B2(KEYINPUT39), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n665), .A2(new_n272), .A3(new_n719), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n894), .B1(new_n915), .B2(new_n923), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n738), .B(new_n465), .C1(KEYINPUT29), .C2(new_n744), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n674), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n770), .A2(new_n765), .A3(new_n767), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n465), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT113), .Z(new_n945));
  AOI21_X1  g0745(.A(new_n874), .B1(new_n917), .B2(new_n919), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n926), .A2(new_n912), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n943), .A2(new_n946), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n934), .A2(new_n933), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n925), .B1(new_n952), .B2(new_n930), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n953), .B2(new_n912), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n954), .B2(new_n949), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n945), .A2(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(G330), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n942), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(KEYINPUT114), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(KEYINPUT114), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n942), .A2(new_n959), .B1(new_n209), .B2(new_n779), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT35), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n510), .A2(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n638), .B(new_n227), .C1(new_n510), .C2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n968), .B2(KEYINPUT110), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(KEYINPUT110), .B2(new_n968), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT36), .Z(new_n971));
  INV_X1    g0771(.A(new_n229), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(G77), .C1(new_n217), .C2(new_n398), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n201), .A2(G68), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n209), .B(G13), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n964), .A2(new_n971), .A3(new_n975), .ZN(G367));
  INV_X1    g0776(.A(new_n784), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n239), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n794), .B1(new_n213), .B2(new_n368), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n782), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n819), .A2(new_n217), .B1(new_n814), .B2(new_n250), .ZN(new_n981));
  INV_X1    g0781(.A(G137), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n286), .B1(new_n807), .B2(new_n982), .C1(new_n398), .C2(new_n810), .ZN(new_n983));
  INV_X1    g0783(.A(new_n862), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n981), .B(new_n983), .C1(new_n801), .C2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n201), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G159), .A2(new_n804), .B1(new_n799), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(new_n860), .C2(new_n825), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n811), .A2(G116), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT46), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT117), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G283), .B2(new_n799), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n819), .A2(new_n206), .B1(new_n814), .B2(new_n205), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n403), .B1(new_n995), .B2(new_n807), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n990), .C2(new_n989), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n804), .A2(G294), .B1(new_n801), .B2(G311), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n825), .A2(new_n632), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n988), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n793), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n678), .A2(new_n707), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(new_n681), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n742), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n844), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT43), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n685), .B(new_n686), .C1(new_n531), .C2(new_n719), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n626), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n686), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(KEYINPUT115), .B(new_n686), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n719), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n690), .A2(new_n707), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT42), .B1(new_n1022), .B2(new_n721), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT42), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n721), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1011), .B(new_n1012), .C1(new_n1020), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1030), .A2(new_n1010), .A3(new_n1009), .A4(new_n1019), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n718), .A2(new_n1022), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT116), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT45), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n721), .A2(new_n722), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n1022), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n723), .A2(new_n1024), .A3(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1022), .A2(KEYINPUT44), .A3(new_n1043), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT44), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n723), .B2(new_n1024), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n717), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1046), .A2(new_n1050), .A3(new_n718), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n720), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n711), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n721), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(new_n716), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n777), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n726), .B(KEYINPUT41), .Z(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n781), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1008), .B1(new_n1041), .B2(new_n1062), .ZN(G387));
  INV_X1    g0863(.A(new_n776), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n775), .B1(new_n745), .B2(new_n772), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n1058), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1058), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n777), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n726), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n794), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n236), .A2(new_n785), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1072), .A2(new_n977), .B1(new_n728), .B2(new_n788), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n366), .A2(new_n337), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT50), .Z(new_n1075));
  AOI21_X1  g0875(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n728), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1073), .A2(new_n1077), .B1(new_n206), .B2(new_n725), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n632), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n804), .B1(new_n799), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n840), .B2(new_n802), .C1(new_n825), .C2(new_n995), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n827), .A2(G283), .B1(new_n811), .B2(G294), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT49), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n419), .B1(G326), .B2(new_n832), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n638), .B2(new_n814), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n807), .A2(new_n860), .B1(new_n810), .B2(new_n250), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT118), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n419), .B1(new_n205), .B2(new_n814), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT119), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n804), .A2(new_n332), .B1(new_n801), .B2(G159), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n577), .A2(new_n827), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n217), .C2(new_n800), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n825), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(G50), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1091), .A2(new_n1092), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n793), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n782), .B1(new_n1071), .B2(new_n1078), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n711), .B2(new_n792), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n781), .B2(new_n1068), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1070), .A2(new_n1107), .ZN(G393));
  AND3_X1   g0908(.A1(new_n1046), .A2(new_n718), .A3(new_n1050), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n718), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n781), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1071), .B1(G97), .B2(new_n725), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n977), .A2(new_n243), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n783), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n825), .A2(new_n808), .B1(new_n860), .B2(new_n802), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT120), .Z(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n819), .A2(new_n250), .B1(new_n814), .B2(new_n425), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G68), .B2(new_n811), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n804), .A2(new_n986), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n799), .A2(new_n366), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n403), .B1(new_n832), .B2(new_n984), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n816), .B(new_n280), .C1(new_n840), .C2(new_n807), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n804), .A2(new_n1079), .B1(G116), .B2(new_n827), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n610), .B2(new_n800), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT121), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1128), .B(new_n1131), .C1(G283), .C2(new_n811), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n825), .A2(new_n829), .B1(new_n995), .B2(new_n802), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT52), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1126), .A2(new_n1127), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1116), .B1(new_n1135), .B2(new_n1104), .C1(new_n1024), .C2(new_n844), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1069), .A2(new_n1054), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n726), .B1(new_n1069), .B2(new_n1054), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1112), .B(new_n1136), .C1(new_n1138), .C2(new_n1139), .ZN(G390));
  AOI21_X1  g0940(.A(new_n922), .B1(new_n694), .B2(new_n882), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n920), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n938), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT39), .B1(new_n953), .B2(new_n912), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n938), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n953), .B2(new_n912), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n732), .B1(new_n541), .B2(new_n684), .ZN(new_n1149));
  AND4_X1   g0949(.A1(new_n692), .A2(new_n537), .A3(new_n540), .A4(new_n581), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n692), .B1(new_n690), .B2(new_n691), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n707), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n922), .B1(new_n1153), .B2(new_n872), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1148), .B1(new_n1154), .B2(new_n1142), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n771), .A2(G330), .A3(new_n875), .A4(new_n920), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1146), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n943), .A2(G330), .A3(new_n946), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n770), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n765), .A2(new_n767), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n875), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1142), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1154), .A2(new_n1156), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n771), .A2(G330), .A3(new_n875), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1158), .B1(new_n1167), .B2(new_n1142), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n1141), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n465), .A2(G330), .A3(new_n943), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n940), .A2(new_n674), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n727), .B1(new_n1161), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT122), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n1172), .C1(new_n1157), .C2(new_n1160), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n883), .A2(new_n873), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1147), .B1(new_n1179), .B2(new_n920), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1155), .B(new_n1156), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n872), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n707), .B(new_n1182), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n920), .B1(new_n1183), .B2(new_n922), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n937), .A2(new_n1143), .B1(new_n1184), .B2(new_n1148), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1181), .B1(new_n1185), .B2(new_n1159), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1175), .B1(new_n1186), .B2(new_n1172), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1174), .B1(new_n1177), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1161), .A2(new_n781), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n877), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n782), .B1(new_n1190), .B2(new_n332), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n280), .B1(new_n832), .B2(G125), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n201), .B2(new_n814), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n811), .A2(G150), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT53), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G159), .C2(new_n827), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT54), .B(G143), .ZN(new_n1197));
  INV_X1    g0997(.A(G128), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n800), .A2(new_n1197), .B1(new_n802), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G137), .B2(new_n804), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1196), .B(new_n1200), .C1(new_n856), .C2(new_n825), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n819), .A2(new_n250), .B1(new_n814), .B2(new_n217), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n812), .B(new_n280), .C1(new_n610), .C2(new_n807), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G97), .C2(new_n799), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n804), .A2(G107), .B1(new_n801), .B2(G283), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n638), .C2(new_n825), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1191), .B1(new_n1207), .B2(new_n793), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1178), .B2(new_n791), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1189), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1188), .A2(new_n1211), .ZN(G378));
  NAND3_X1  g1012(.A1(new_n378), .A2(new_n355), .A3(new_n382), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n893), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(new_n379), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n955), .A2(G330), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n955), .B2(G330), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n939), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n953), .A2(new_n912), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n949), .B1(new_n1226), .B2(new_n947), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n915), .A2(KEYINPUT40), .A3(new_n951), .ZN(new_n1228));
  OAI21_X1  g1028(.A(G330), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1221), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n894), .B1(new_n923), .B2(new_n915), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1147), .B2(new_n1178), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n955), .A2(G330), .A3(new_n1222), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1225), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1171), .B1(new_n1186), .B2(new_n1172), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(KEYINPUT57), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1160), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1173), .A2(new_n1238), .A3(new_n1181), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1239), .A2(new_n1171), .B1(new_n1225), .B2(new_n1234), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1237), .B(new_n726), .C1(new_n1240), .C2(KEYINPUT57), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1222), .A2(new_n791), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n782), .B1(new_n1190), .B2(new_n986), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1101), .A2(G107), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n403), .A2(new_n300), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n819), .A2(new_n217), .B1(new_n807), .B2(new_n834), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n810), .A2(new_n250), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n814), .A2(new_n398), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n801), .A2(G116), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n577), .A2(new_n799), .B1(new_n804), .B2(G97), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1244), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT58), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G50), .B1(new_n278), .B2(new_n300), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1252), .A2(new_n1253), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G132), .A2(new_n804), .B1(new_n799), .B2(G137), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n801), .A2(G125), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1197), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n827), .A2(G150), .B1(new_n811), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G128), .B2(new_n1101), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n815), .A2(G159), .ZN(new_n1264));
  AOI211_X1 g1064(.A(G33), .B(G41), .C1(new_n832), .C2(G124), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1255), .B1(new_n1253), .B2(new_n1252), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1243), .B1(new_n1268), .B2(new_n793), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1235), .A2(new_n781), .B1(new_n1242), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1241), .A2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n1169), .A2(new_n781), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n782), .B1(new_n1190), .B2(G68), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n206), .A2(new_n800), .B1(new_n861), .B2(new_n638), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G294), .B2(new_n801), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1101), .A2(G283), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n280), .B1(new_n807), .B2(new_n835), .C1(new_n250), .C2(new_n814), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G97), .B2(new_n811), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1275), .A2(new_n1099), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1248), .B1(G159), .B2(new_n811), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n337), .B2(new_n819), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n403), .B(new_n1281), .C1(G128), .C2(new_n832), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n860), .B2(new_n800), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n804), .A2(new_n1258), .B1(new_n801), .B2(G132), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n825), .B2(new_n982), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT123), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1279), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1273), .B1(new_n1287), .B2(new_n793), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n790), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n920), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1272), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1172), .A2(new_n1061), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(G381));
  NAND2_X1  g1095(.A1(new_n1112), .A2(new_n1136), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1139), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1137), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n891), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1070), .A2(new_n848), .A3(new_n1107), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1300), .A2(G381), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(G378), .A2(new_n1299), .A3(new_n1301), .A4(G387), .ZN(new_n1302));
  INV_X1    g1102(.A(G375), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G407));
  AOI21_X1  g1104(.A(new_n701), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n701), .A2(G343), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(G378), .A2(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1303), .A2(KEYINPUT124), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT124), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1305), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1305), .B(KEYINPUT125), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G409));
  NAND3_X1  g1115(.A1(new_n1241), .A2(G378), .A3(new_n1270), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT122), .B1(new_n1161), .B2(new_n1173), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1176), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1210), .B1(new_n1318), .B2(new_n1174), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1235), .A2(new_n1236), .A3(new_n1061), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1270), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1306), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT60), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1324), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n727), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1167), .A2(new_n1142), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1159), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1179), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n940), .A2(new_n674), .A3(new_n1170), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(KEYINPUT60), .A3(new_n1330), .A4(new_n1166), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1325), .A2(new_n1326), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(KEYINPUT126), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1325), .A2(new_n1326), .A3(new_n1331), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1292), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n891), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(G384), .A3(new_n1292), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1306), .A2(G2897), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1340), .ZN(new_n1342));
  AOI21_X1  g1142(.A(G384), .B1(new_n1336), .B2(new_n1292), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n891), .B(new_n1291), .C1(new_n1333), .C2(new_n1335), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(KEYINPUT63), .B1(new_n1323), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1323), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G387), .A2(new_n1298), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1066), .B1(new_n1068), .B2(new_n1111), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n780), .B1(new_n1352), .B2(new_n1060), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1037), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1354));
  AOI211_X1 g1154(.A(new_n1034), .B(new_n1033), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1357), .A2(G390), .A3(new_n1008), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1300), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n848), .B1(new_n1070), .B2(new_n1107), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1351), .A2(new_n1358), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1361), .B1(new_n1351), .B2(new_n1358), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1362), .A2(new_n1363), .A3(KEYINPUT61), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1365), .A2(new_n1348), .A3(KEYINPUT63), .A4(new_n1307), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1350), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1323), .A2(new_n1369), .A3(new_n1348), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT61), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1371), .B1(new_n1323), .B2(new_n1346), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1369), .B1(new_n1323), .B2(new_n1348), .ZN(new_n1373));
  NOR3_X1   g1173(.A1(new_n1370), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT127), .ZN(new_n1375));
  NOR3_X1   g1175(.A1(new_n1362), .A2(new_n1363), .A3(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1351), .A2(new_n1358), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1361), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1351), .A2(new_n1358), .A3(new_n1361), .ZN(new_n1380));
  AOI21_X1  g1180(.A(KEYINPUT127), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1376), .A2(new_n1381), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1368), .B1(new_n1374), .B2(new_n1382), .ZN(G405));
  NAND2_X1  g1183(.A1(G375), .A2(new_n1319), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1384), .A2(new_n1316), .ZN(new_n1385));
  OAI21_X1  g1185(.A(new_n1375), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1379), .A2(KEYINPUT127), .A3(new_n1380), .ZN(new_n1387));
  INV_X1    g1187(.A(new_n1348), .ZN(new_n1388));
  AND3_X1   g1188(.A1(new_n1386), .A2(new_n1387), .A3(new_n1388), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1388), .B1(new_n1386), .B2(new_n1387), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1385), .B1(new_n1389), .B2(new_n1390), .ZN(new_n1391));
  OAI21_X1  g1191(.A(new_n1348), .B1(new_n1376), .B2(new_n1381), .ZN(new_n1392));
  INV_X1    g1192(.A(new_n1385), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1386), .A2(new_n1387), .A3(new_n1388), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1392), .A2(new_n1393), .A3(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1391), .A2(new_n1395), .ZN(G402));
endmodule


