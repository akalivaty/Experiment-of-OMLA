//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT66), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(G137), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n461), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n472), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n471), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n466), .A2(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n464), .A2(new_n479), .A3(new_n465), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G124), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT68), .Z(G162));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n474), .B2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n474), .A2(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(new_n465), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n481), .A2(G102), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT4), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n464), .A2(G138), .A3(new_n471), .A4(new_n465), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n512), .A2(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT70), .B(G51), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT71), .B(G89), .ZN(new_n531));
  OAI221_X1 g106(.A(new_n529), .B1(new_n519), .B2(new_n530), .C1(new_n517), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n517), .A2(new_n539), .B1(new_n519), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n509), .A2(new_n511), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n517), .A2(new_n549), .B1(new_n519), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n544), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT74), .Z(new_n564));
  XNOR2_X1  g139(.A(new_n517), .B(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G91), .ZN(new_n566));
  INV_X1    g141(.A(new_n519), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G53), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n565), .A2(G87), .ZN(new_n573));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n514), .B1(new_n544), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n567), .B2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G288));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n512), .A2(new_n578), .A3(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT75), .B1(new_n544), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G48), .B2(new_n567), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n586));
  OAI21_X1  g161(.A(G86), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G305));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n517), .A2(new_n589), .B1(new_n519), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n514), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n544), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(G54), .A2(new_n567), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n565), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n565), .B2(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  XOR2_X1   g185(.A(G299), .B(KEYINPUT77), .Z(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G860), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n606), .B1(G559), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT78), .Z(G148));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n552), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n606), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n489), .A2(G123), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n479), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n486), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G135), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2100), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(G2451), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n645), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n651), .A4(new_n643), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n646), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n638), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  INV_X1    g231(.A(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n658), .B2(new_n637), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n668), .A2(KEYINPUT17), .A3(new_n665), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n668), .B2(KEYINPUT17), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n669), .A2(new_n670), .A3(new_n664), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n681), .B2(new_n683), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1991), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n680), .A2(new_n683), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n690), .A2(new_n691), .A3(new_n687), .A4(new_n684), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G1991), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n694), .A3(G1996), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(G1996), .B1(new_n692), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n694), .ZN(new_n701));
  INV_X1    g276(.A(G1996), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n700), .B1(new_n703), .B2(new_n695), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n676), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n700), .A3(new_n695), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n707), .A3(new_n675), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT29), .Z(new_n713));
  INV_X1    g288(.A(G2090), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G4), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n607), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT89), .B(G1348), .Z(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n710), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n466), .A2(G140), .A3(new_n467), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n489), .A2(G128), .ZN(new_n725));
  OAI221_X1 g300(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n471), .C2(G116), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT91), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT93), .B(G2067), .Z(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NOR4_X1   g309(.A1(new_n715), .A2(new_n720), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT24), .B(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(new_n710), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT97), .Z(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n483), .B2(new_n710), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(G16), .ZN(new_n742));
  MUX2_X1   g317(.A(G19), .B(new_n552), .S(new_n742), .Z(new_n743));
  XOR2_X1   g318(.A(KEYINPUT90), .B(G1341), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n741), .B(new_n745), .C1(G29), .C2(new_n630), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT31), .B(G11), .Z(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n710), .B1(new_n748), .B2(G28), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(new_n750), .B1(new_n748), .B2(G28), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(G171), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G5), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n716), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n716), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n756), .C2(new_n755), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(G1966), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n628), .A2(G141), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n489), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n767), .A2(new_n768), .B1(G105), .B2(new_n481), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G32), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n762), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n746), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G20), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n742), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  INV_X1    g355(.A(G299), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n716), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(G29), .A2(G33), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT96), .B1(new_n486), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT25), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n476), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n788), .A2(new_n789), .B1(new_n479), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n786), .B(new_n793), .C1(new_n789), .C2(new_n788), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n486), .A2(KEYINPUT96), .A3(new_n785), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n784), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2072), .ZN(new_n798));
  NOR2_X1   g373(.A1(G27), .A2(G29), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G164), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(G2078), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n777), .A2(new_n783), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n713), .A2(new_n714), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n735), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G22), .B(G303), .S(new_n742), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT88), .B(G1971), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G288), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G16), .B2(G23), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n716), .A2(G6), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G305), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT87), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n710), .A2(G25), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n628), .A2(KEYINPUT85), .A3(G131), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT85), .ZN(new_n826));
  INV_X1    g401(.A(G131), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n486), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n489), .A2(G119), .ZN(new_n830));
  OAI221_X1 g405(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n471), .C2(G107), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n824), .B1(new_n833), .B2(G29), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT35), .B(G1991), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  MUX2_X1   g412(.A(G24), .B(G290), .S(new_n742), .Z(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1986), .Z(new_n839));
  OR2_X1    g414(.A1(new_n834), .A2(new_n836), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n823), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n805), .B1(new_n842), .B2(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(new_n805), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(G150));
  INV_X1    g422(.A(new_n517), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n848), .A2(G93), .B1(G55), .B2(new_n567), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n514), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n607), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n851), .B(new_n552), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT100), .Z(new_n861));
  OAI21_X1  g436(.A(new_n614), .B1(new_n859), .B2(KEYINPUT39), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(G145));
  XOR2_X1   g438(.A(new_n483), .B(KEYINPUT102), .Z(new_n864));
  XOR2_X1   g439(.A(G162), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT103), .A3(G142), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  INV_X1    g444(.A(G142), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n486), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n489), .A2(G130), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT104), .ZN(new_n874));
  OAI221_X1 g449(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n471), .C2(G118), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n633), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n829), .A2(new_n877), .A3(new_n832), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n829), .B2(new_n832), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n876), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n867), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n884), .A3(new_n867), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n730), .A2(new_n796), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n728), .B(new_n729), .C1(new_n794), .C2(new_n795), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n503), .A2(new_n504), .ZN(new_n891));
  INV_X1    g466(.A(new_n501), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n506), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n499), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n770), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n890), .A2(new_n896), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n886), .A2(new_n887), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n890), .A2(new_n896), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n885), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n899), .A2(new_n902), .A3(new_n630), .ZN(new_n903));
  INV_X1    g478(.A(new_n630), .ZN(new_n904));
  INV_X1    g479(.A(new_n887), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n905), .A2(new_n885), .B1(new_n900), .B2(new_n901), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n886), .A2(new_n897), .A3(new_n898), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n866), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n630), .B1(new_n899), .B2(new_n902), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n904), .A3(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n865), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(G395));
  NAND2_X1  g491(.A1(new_n851), .A2(new_n617), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n606), .A2(new_n781), .ZN(new_n918));
  OAI211_X1 g493(.A(G299), .B(new_n601), .C1(new_n605), .C2(new_n604), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n919), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n606), .A2(new_n781), .A3(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n921), .A2(new_n922), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n619), .B(new_n857), .ZN(new_n933));
  MUX2_X1   g508(.A(new_n920), .B(new_n932), .S(new_n933), .Z(new_n934));
  XNOR2_X1  g509(.A(G166), .B(G305), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n809), .A2(G290), .ZN(new_n936));
  AOI21_X1  g511(.A(G288), .B1(new_n595), .B2(new_n593), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n934), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n917), .B1(new_n943), .B2(new_n617), .ZN(G295));
  OAI21_X1  g519(.A(new_n917), .B1(new_n943), .B2(new_n617), .ZN(G331));
  INV_X1    g520(.A(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(G286), .A2(G301), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n534), .B2(new_n535), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n857), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(G168), .A2(G171), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n858), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n953), .B(new_n930), .C1(new_n923), .C2(new_n928), .ZN(new_n954));
  INV_X1    g529(.A(new_n953), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n920), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n946), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n929), .A2(new_n931), .A3(new_n955), .ZN(new_n958));
  INV_X1    g533(.A(new_n956), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n940), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n913), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n950), .A2(new_n952), .A3(KEYINPUT41), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n940), .B1(new_n920), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n955), .A2(KEYINPUT41), .A3(new_n927), .A4(new_n925), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n960), .A2(new_n967), .A3(new_n962), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(KEYINPUT44), .B2(new_n972), .ZN(G397));
  AOI21_X1  g548(.A(G1384), .B1(new_n893), .B2(new_n894), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT112), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n730), .B(G2067), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(G1996), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n771), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n979), .A2(new_n980), .B1(KEYINPUT111), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n770), .ZN(new_n984));
  OAI221_X1 g559(.A(new_n983), .B1(KEYINPUT111), .B2(new_n982), .C1(new_n702), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n833), .A2(new_n835), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n829), .A2(new_n836), .A3(new_n832), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n991));
  INV_X1    g566(.A(new_n978), .ZN(new_n992));
  AND2_X1   g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n502), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT69), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n501), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n998), .B(new_n999), .C1(new_n1002), .C2(new_n499), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT50), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n977), .B1(new_n974), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1004), .A2(G2084), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n997), .A2(new_n1008), .A3(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n976), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1966), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(G8), .B(G286), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1007), .A2(new_n1011), .A3(G286), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT123), .B(new_n1013), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n998), .B1(new_n895), .B2(new_n999), .ZN(new_n1017));
  NOR3_X1   g592(.A1(G164), .A2(KEYINPUT115), .A3(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1005), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1006), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n740), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(G168), .C1(G1966), .C2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT123), .B1(new_n1026), .B2(new_n1013), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1012), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n1012), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(new_n1008), .C1(G164), .C2(G1384), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1010), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1036), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n714), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT55), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(G8), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n997), .A2(new_n1003), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1015), .B1(new_n1048), .B2(new_n977), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n809), .A2(G1976), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT116), .B(G1981), .Z(new_n1054));
  NAND3_X1  g629(.A1(new_n584), .A2(new_n587), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT117), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n584), .A2(new_n587), .A3(new_n1057), .A4(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT118), .B(G86), .Z(new_n1060));
  OAI21_X1  g635(.A(new_n584), .B1(new_n517), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1049), .A3(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1053), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1037), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n997), .A2(KEYINPUT50), .A3(new_n1003), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n976), .B1(new_n974), .B2(new_n1005), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G2090), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1045), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1047), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1035), .B2(G2078), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1961), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT45), .B(new_n999), .C1(new_n1002), .C2(new_n499), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n977), .A3(KEYINPUT53), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1008), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT124), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n756), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1048), .A2(KEYINPUT45), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1090), .B(new_n1091), .C1(new_n1092), .C2(new_n1086), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1082), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1079), .A2(G301), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1029), .A2(new_n1031), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1067), .A2(new_n1051), .A3(new_n809), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1059), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1049), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1047), .B2(new_n1070), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  OAI211_X1 g676(.A(G8), .B(G168), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1079), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1043), .A2(G8), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1045), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1101), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1047), .A3(new_n1071), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1096), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G171), .B(KEYINPUT54), .ZN(new_n1110));
  INV_X1    g685(.A(new_n975), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(new_n1010), .A3(KEYINPUT53), .A4(new_n1085), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1081), .A2(new_n1090), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1094), .B2(new_n1110), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1079), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1028), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1032), .A2(new_n1010), .A3(new_n702), .A4(new_n1034), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1048), .A2(new_n977), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n553), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT59), .B(new_n553), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT120), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1032), .A2(new_n1010), .A3(new_n1034), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT119), .B(G1956), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G299), .B(KEYINPUT57), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1137), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1075), .A2(new_n1134), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n1132), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1129), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1139), .A3(new_n1132), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT61), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1127), .A2(new_n1128), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT61), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT61), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(KEYINPUT122), .A3(new_n1128), .A4(new_n1127), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1120), .A2(G2067), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1041), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n719), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(KEYINPUT60), .B2(new_n607), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1148), .A2(new_n1152), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1143), .B1(new_n1155), .B2(new_n606), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1144), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1116), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n996), .B1(new_n1109), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n981), .B(KEYINPUT46), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n979), .A2(new_n980), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n984), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT47), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n991), .B(KEYINPUT48), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n990), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n985), .A2(new_n987), .B1(G2067), .B2(new_n730), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n979), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1163), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(G227), .A2(new_n458), .ZN(new_n1174));
  NAND4_X1  g748(.A1(new_n705), .A2(new_n660), .A3(new_n708), .A4(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g749(.A(new_n1175), .B(KEYINPUT126), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n914), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g751(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n972), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n1179));
  INV_X1    g753(.A(new_n971), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NAND4_X1  g756(.A1(new_n1181), .A2(new_n1182), .A3(new_n914), .A4(new_n1176), .ZN(new_n1183));
  AND2_X1   g757(.A1(new_n1178), .A2(new_n1183), .ZN(G308));
  NAND2_X1  g758(.A1(new_n1178), .A2(new_n1183), .ZN(G225));
endmodule


