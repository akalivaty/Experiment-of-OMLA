//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT68), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n473), .A2(new_n474), .A3(new_n477), .A4(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n469), .B1(new_n480), .B2(G2105), .ZN(G160));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(new_n464), .B2(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT71), .Z(new_n485));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  AOI22_X1  g061(.A1(G136), .A2(new_n466), .B1(new_n486), .B2(G2104), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n482), .A2(G102), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n482), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n491), .A2(G2104), .B1(G126), .B2(new_n483), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n482), .A2(G138), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n473), .A3(new_n474), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n482), .C1(new_n471), .C2(new_n472), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT74), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(G50), .A2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n518), .A2(G651), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NOR2_X1   g097(.A1(new_n508), .A2(KEYINPUT76), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n511), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(G543), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n514), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n505), .A2(KEYINPUT75), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT75), .B1(new_n505), .B2(new_n530), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n509), .A2(new_n513), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT77), .B(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI221_X1 g118(.A(new_n540), .B1(new_n541), .B2(new_n542), .C1(new_n526), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n527), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n514), .A2(G81), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n539), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT79), .Z(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n523), .C2(new_n525), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n505), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n514), .A2(G91), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  AND2_X1   g143(.A1(new_n546), .A2(new_n547), .ZN(G301));
  NAND2_X1  g144(.A1(new_n514), .A2(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(G49), .B(G543), .C1(new_n523), .C2(new_n525), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n505), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(G651), .B1(new_n511), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n509), .A2(G86), .A3(new_n513), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n539), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n541), .B2(new_n583), .C1(new_n526), .C2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G171), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n526), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(G54), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n509), .A2(G92), .A3(new_n513), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n539), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT81), .B1(new_n602), .B2(new_n590), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n593), .B1(new_n591), .B2(new_n603), .ZN(G284));
  OAI21_X1  g179(.A(new_n593), .B1(new_n591), .B2(new_n603), .ZN(G321));
  NOR2_X1   g180(.A1(G286), .A2(new_n590), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n590), .ZN(G297));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n590), .ZN(G280));
  INV_X1    g184(.A(new_n602), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n553), .A2(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n602), .A2(G559), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g191(.A1(new_n473), .A2(new_n474), .A3(new_n467), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n619), .B2(new_n618), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n620), .A3(new_n621), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n466), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(G111), .A2(G2105), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G99), .B2(new_n482), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n463), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2427), .ZN(new_n639));
  INV_X1    g214(.A(G2430), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  INV_X1    g234(.A(new_n655), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n662), .B2(new_n653), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n654), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n654), .A2(new_n657), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n660), .B1(new_n665), .B2(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n659), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n632), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n621), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n675), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT20), .Z(new_n679));
  AOI211_X1 g254(.A(new_n677), .B(new_n679), .C1(new_n672), .C2(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  NAND3_X1  g263(.A1(new_n587), .A2(G16), .A3(new_n588), .ZN(new_n689));
  OR2_X1    g264(.A1(G16), .A2(G24), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(KEYINPUT89), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1986), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n697), .A3(new_n694), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G166), .A2(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G16), .B2(G22), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(G1971), .C1(G16), .C2(G22), .ZN(new_n704));
  INV_X1    g279(.A(G305), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G6), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n703), .B(new_n704), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  OAI21_X1  g293(.A(KEYINPUT34), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n703), .A2(new_n704), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n716), .B(new_n717), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n710), .A2(new_n711), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n466), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n483), .A2(G119), .ZN(new_n726));
  AND2_X1   g301(.A1(G107), .A2(G2105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G95), .B2(new_n482), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n726), .C1(new_n463), .C2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT87), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT87), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G25), .B(new_n729), .S(new_n734), .Z(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT88), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n719), .A2(new_n724), .A3(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(KEYINPUT90), .B(KEYINPUT36), .C1(new_n699), .C2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n724), .A2(new_n738), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n696), .A2(new_n698), .ZN(new_n742));
  NAND2_X1  g317(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n719), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n466), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n467), .A2(G105), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n730), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n730), .B2(G32), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  INV_X1    g333(.A(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n759), .B2(KEYINPUT30), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n762), .A2(new_n759), .A3(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n759), .B2(KEYINPUT30), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n758), .B1(new_n761), .B2(new_n766), .C1(new_n631), .C2(new_n733), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n756), .A2(new_n757), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n730), .A2(G33), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n467), .A2(G103), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT92), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n466), .A2(G139), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n473), .A2(new_n474), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n774), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n773), .C1(new_n482), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G1966), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n713), .A2(G21), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G286), .B2(G16), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n768), .B(new_n779), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n554), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n733), .A2(G26), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT28), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n787), .B(KEYINPUT91), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G128), .ZN(new_n794));
  MUX2_X1   g369(.A(G104), .B(G116), .S(G2105), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2104), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G140), .B2(new_n466), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n790), .B(new_n793), .C1(new_n730), .C2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G164), .A2(new_n734), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G27), .B2(new_n734), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n783), .A2(new_n786), .A3(new_n807), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n777), .A2(KEYINPUT93), .A3(new_n778), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT93), .B1(new_n777), .B2(new_n778), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G34), .ZN(new_n811));
  AOI22_X1  g386(.A1(G160), .A2(G29), .B1(new_n733), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n809), .A2(new_n810), .B1(G2084), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G4), .A2(G16), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n610), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n733), .A2(G35), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G162), .B2(new_n733), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT100), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n808), .A2(new_n813), .A3(new_n817), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n713), .A2(G5), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G171), .B2(new_n713), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(KEYINPUT97), .B(new_n828), .C1(G171), .C2(new_n713), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1961), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n822), .A2(KEYINPUT100), .A3(new_n823), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n782), .A2(new_n780), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT96), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n812), .A2(G2084), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT98), .Z(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n713), .A2(G20), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G299), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1956), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n835), .A2(new_n837), .A3(new_n839), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n827), .A2(new_n834), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n745), .A2(KEYINPUT102), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT102), .B1(new_n745), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n745), .A2(new_n846), .ZN(G150));
  AOI22_X1  g425(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n539), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n514), .B2(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(new_n526), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT103), .B(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n553), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n610), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n858), .B1(new_n866), .B2(new_n867), .ZN(G145));
  NAND2_X1  g443(.A1(new_n483), .A2(G130), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT106), .B1(new_n482), .B2(G118), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n482), .A2(KEYINPUT106), .A3(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n466), .ZN(new_n874));
  INV_X1    g449(.A(G142), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n874), .A2(KEYINPUT105), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT105), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(new_n618), .Z(new_n879));
  XOR2_X1   g454(.A(new_n729), .B(KEYINPUT107), .Z(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n798), .B(new_n501), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n776), .B(new_n751), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g465(.A(G160), .B(new_n631), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g473(.A1(new_n855), .A2(new_n590), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n614), .B(new_n859), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n610), .A2(new_n607), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n602), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n901), .A2(new_n906), .A3(KEYINPUT108), .A4(new_n907), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n901), .A2(new_n904), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G290), .A2(G288), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n587), .A2(new_n715), .A3(new_n588), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G303), .B(new_n705), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n900), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n912), .A2(new_n911), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n924), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n910), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n913), .A2(new_n925), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n899), .B1(new_n931), .B2(new_n590), .ZN(G295));
  OAI21_X1  g507(.A(new_n899), .B1(new_n931), .B2(new_n590), .ZN(G331));
  XNOR2_X1  g508(.A(new_n554), .B(new_n855), .ZN(new_n934));
  AOI21_X1  g509(.A(G286), .B1(new_n546), .B2(new_n547), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n546), .A2(G286), .A3(new_n547), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n939), .A2(new_n859), .A3(new_n935), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n906), .B(new_n907), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n859), .B1(new_n939), .B2(new_n935), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n934), .A3(new_n937), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n903), .A4(new_n902), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n921), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n895), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n921), .B1(new_n941), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n895), .A4(new_n945), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n948), .B2(new_n951), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(G397));
  AOI21_X1  g530(.A(G1384), .B1(new_n492), .B2(new_n500), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n478), .A2(new_n479), .ZN(new_n959));
  OAI21_X1  g534(.A(G2105), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(G40), .A3(new_n468), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(new_n752), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT110), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n798), .B(G2067), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n963), .B2(new_n752), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n737), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n729), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n729), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(G290), .B(G1986), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n962), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n961), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n497), .A2(new_n499), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n483), .A2(G126), .ZN(new_n980));
  INV_X1    g555(.A(new_n489), .ZN(new_n981));
  INV_X1    g556(.A(G114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT72), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT72), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G114), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n986), .B2(G2105), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n980), .B1(new_n987), .B2(new_n463), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n978), .C1(new_n979), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n956), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n977), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n995));
  NAND3_X1  g570(.A1(new_n501), .A2(new_n978), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(new_n956), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n998), .A2(G2084), .A3(new_n961), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(G286), .C1(new_n994), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT122), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1003), .B(new_n469), .C1(new_n480), .C2(G2105), .ZN(new_n1004));
  AND4_X1   g579(.A1(KEYINPUT117), .A2(new_n501), .A3(KEYINPUT45), .A4(new_n978), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT117), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n957), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n780), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n998), .A2(new_n961), .ZN(new_n1009));
  INV_X1    g584(.A(G2084), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(KEYINPUT122), .A3(G8), .A4(G286), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(G8), .C1(new_n1012), .C2(G286), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G286), .A2(G8), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n780), .A2(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT51), .B(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT62), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT62), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G160), .A2(G40), .A3(new_n956), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n570), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n578), .A2(new_n579), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n578), .B2(new_n579), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT113), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT113), .B(new_n1035), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(G8), .A3(new_n1026), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(G8), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1029), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n989), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n956), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n957), .A2(new_n1004), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n702), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1009), .A2(new_n823), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1019), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1041), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n956), .A2(new_n997), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n956), .A2(new_n1055), .A3(new_n997), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n956), .A2(new_n995), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n961), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n823), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1046), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT116), .A3(new_n1050), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n977), .A2(new_n993), .A3(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT123), .B(G1961), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n998), .B2(new_n961), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1045), .B2(G2078), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1019), .B1(new_n1046), .B2(new_n1060), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1051), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n1052), .A2(new_n1063), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1022), .A2(new_n1025), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1026), .A2(G8), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1037), .A2(new_n1038), .A3(new_n715), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1031), .B(KEYINPUT114), .Z(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1041), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1084));
  INV_X1    g659(.A(G1956), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n563), .A2(new_n567), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(G299), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT56), .B(G2072), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n977), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n816), .B1(new_n998), .B2(new_n961), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1004), .A2(new_n800), .A3(new_n956), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n602), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(new_n1089), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1045), .A2(new_n1092), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1956), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1096), .A2(new_n602), .A3(new_n1097), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT60), .B1(new_n1105), .B2(new_n1098), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n610), .A2(new_n1096), .A3(new_n1107), .A4(new_n1097), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT120), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1026), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1045), .B2(G1996), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n554), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1112), .B2(new_n554), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1106), .B(new_n1108), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT61), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1103), .A2(KEYINPUT61), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1104), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G301), .B(KEYINPUT54), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1070), .A3(new_n1069), .ZN(new_n1125));
  AND4_X1   g700(.A1(G40), .A2(new_n957), .A3(new_n468), .A4(new_n1065), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n480), .B(KEYINPUT124), .Z(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n1091), .C1(new_n482), .C2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1128), .A2(new_n1070), .A3(new_n1068), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1063), .A2(new_n1052), .A3(new_n1074), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1023), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1076), .B(new_n1083), .C1(new_n1123), .C2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1018), .A2(new_n1019), .A3(G286), .ZN(new_n1136));
  AND4_X1   g711(.A1(KEYINPUT63), .A2(new_n1135), .A3(new_n1052), .A4(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1063), .A2(new_n1052), .A3(new_n1074), .A4(new_n1136), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT118), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1137), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n975), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n1146));
  INV_X1    g721(.A(new_n962), .ZN(new_n1147));
  NOR3_X1   g722(.A1(G290), .A2(new_n1147), .A3(G1986), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n973), .B2(KEYINPUT126), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n962), .A2(new_n963), .ZN(new_n1154));
  NOR2_X1   g729(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n966), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n962), .B1(new_n1157), .B2(new_n751), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1156), .B(new_n1158), .C1(new_n1154), .C2(new_n1153), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n968), .A2(new_n971), .B1(new_n800), .B2(new_n798), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1147), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1152), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g739(.A1(new_n948), .A2(new_n951), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G401), .A2(new_n460), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n687), .A2(new_n669), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n897), .A3(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


