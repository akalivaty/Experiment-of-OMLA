//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n468), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(G136), .B2(new_n467), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(new_n490), .A3(new_n486), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n478), .B2(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G166));
  XOR2_X1   g086(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G89), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(new_n506), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n499), .A2(new_n500), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n501), .A2(KEYINPUT70), .A3(G63), .A4(G651), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n520), .A2(new_n521), .B1(G51), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n516), .B1(KEYINPUT71), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n503), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n506), .A2(new_n533), .B1(new_n508), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n503), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n506), .A2(new_n542), .B1(new_n508), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n525), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n503), .ZN(new_n554));
  INV_X1    g129(.A(new_n506), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G91), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n554), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G299));
  INV_X1    g137(.A(new_n538), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n536), .A2(KEYINPUT73), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT75), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n537), .B2(new_n538), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G166), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n525), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n501), .A2(new_n505), .A3(G87), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n499), .B2(new_n500), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n501), .A2(new_n505), .A3(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n525), .A2(G48), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  INV_X1    g156(.A(G72), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n518), .A2(new_n581), .B1(new_n582), .B2(new_n522), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI221_X1 g160(.A(KEYINPUT76), .B1(new_n582), .B2(new_n522), .C1(new_n518), .C2(new_n581), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(G651), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n555), .A2(G85), .B1(G47), .B2(new_n525), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G290));
  AND3_X1   g166(.A1(new_n501), .A2(new_n505), .A3(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G301), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G284));
  AOI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G286), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n561), .B(KEYINPUT78), .Z(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G297));
  AOI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G280));
  INV_X1    g182(.A(new_n598), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n489), .A2(new_n469), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(G2100), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n467), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n468), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n619), .A2(new_n620), .A3(new_n627), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(G401));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n618), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n626), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n658), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n658), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT81), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n671), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G25), .A2(G29), .ZN(new_n682));
  OR2_X1    g257(.A1(G95), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT82), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n467), .A2(G131), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n478), .A2(G119), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n682), .B1(new_n689), .B2(G29), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT35), .B(G1991), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT83), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT85), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n694), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n698), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n709));
  OAI21_X1  g284(.A(new_n693), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G290), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G16), .B2(G24), .ZN(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n710), .B(new_n716), .C1(new_n715), .C2(new_n714), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT36), .Z(new_n718));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G29), .B2(G32), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G129), .B2(new_n478), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT89), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  MUX2_X1   g302(.A(new_n719), .B(new_n720), .S(new_n727), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT91), .Z(new_n731));
  NOR2_X1   g306(.A1(G168), .A2(new_n694), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n694), .B2(G21), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NOR2_X1   g309(.A1(G5), .A2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT92), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G171), .B2(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G1961), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n733), .A2(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n694), .A2(G4), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n608), .B2(new_n694), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT86), .Z(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n740), .B2(new_n739), .C1(new_n744), .C2(G1348), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n694), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n561), .B2(new_n694), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1956), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n744), .A2(G1348), .ZN(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G19), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n545), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT87), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1341), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n731), .A2(new_n745), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n757), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2090), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT94), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(G33), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n489), .A2(G127), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n468), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n765), .B(new_n768), .C1(G139), .C2(new_n467), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n763), .B1(new_n769), .B2(new_n757), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2072), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(G160), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n757), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2084), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT31), .B(G11), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n625), .A2(new_n757), .ZN(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT30), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n778), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  NOR2_X1   g359(.A1(G164), .A2(new_n757), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G27), .B2(new_n757), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n777), .B(new_n783), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n771), .B(new_n787), .C1(new_n784), .C2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n757), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT28), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n467), .A2(G140), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G116), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n478), .B2(G128), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n790), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2067), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n788), .B(new_n800), .C1(G1961), .C2(new_n738), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n760), .A2(G2090), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n728), .A2(new_n729), .B1(new_n734), .B2(new_n733), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n718), .A2(new_n756), .A3(new_n762), .A4(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  AOI22_X1  g381(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n503), .ZN(new_n808));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  INV_X1    g384(.A(G55), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n506), .A2(new_n809), .B1(new_n508), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G860), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT37), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n608), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n545), .A2(new_n812), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n541), .A2(new_n544), .B1(new_n808), .B2(new_n811), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n813), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n815), .B1(new_n823), .B2(new_n824), .ZN(G145));
  AND3_X1   g400(.A1(new_n488), .A2(KEYINPUT96), .A3(new_n491), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT96), .B1(new_n488), .B2(new_n491), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n496), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n798), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n467), .A2(G142), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n478), .A2(G130), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n468), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n688), .B(new_n616), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n726), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n769), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n725), .B2(new_n769), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n837), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(G160), .B(new_n625), .ZN(new_n842));
  XNOR2_X1  g417(.A(G162), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n837), .A2(new_n840), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n837), .A2(new_n840), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g426(.A(G290), .B(G305), .ZN(new_n852));
  XNOR2_X1  g427(.A(G166), .B(new_n704), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT42), .ZN(new_n855));
  INV_X1    g430(.A(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n852), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n611), .B(new_n821), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n608), .B1(new_n559), .B2(new_n560), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n559), .A2(new_n608), .A3(new_n560), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(KEYINPUT41), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n866));
  INV_X1    g441(.A(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n864), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n872), .B2(new_n866), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n861), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n861), .ZN(new_n876));
  INV_X1    g451(.A(new_n872), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n860), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n855), .B(new_n859), .C1(new_n875), .C2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G868), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n812), .A2(G868), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G295));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  AOI211_X1 g463(.A(KEYINPUT98), .B(new_n884), .C1(new_n882), .C2(G868), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G331));
  XOR2_X1   g465(.A(new_n821), .B(KEYINPUT99), .Z(new_n891));
  OAI21_X1  g466(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n537), .A2(new_n566), .A3(new_n538), .ZN(new_n893));
  AOI21_X1  g468(.A(G286), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(G286), .A2(new_n538), .A3(new_n537), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n821), .B(KEYINPUT99), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(new_n895), .C1(G301), .C2(G286), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n872), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n872), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT100), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n871), .B2(new_n874), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n906), .B2(new_n854), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n901), .B1(new_n900), .B2(new_n872), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT97), .B1(new_n865), .B2(new_n868), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n897), .B(new_n899), .C1(new_n909), .C2(new_n873), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n857), .A3(new_n902), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT43), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n857), .B1(new_n911), .B2(new_n902), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n869), .A2(new_n897), .A3(new_n899), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n857), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n869), .A2(new_n897), .A3(new_n899), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n900), .B2(new_n872), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NOR4_X1   g496(.A1(new_n914), .A2(new_n920), .A3(new_n921), .A4(G37), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n913), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n907), .B2(new_n912), .ZN(new_n925));
  NOR4_X1   g500(.A1(new_n914), .A2(new_n920), .A3(KEYINPUT43), .A4(G37), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n828), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n470), .A2(G40), .A3(new_n474), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n725), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT104), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n937), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n838), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n798), .A2(G2067), .ZN(new_n942));
  INV_X1    g517(.A(G2067), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n793), .A2(new_n943), .A3(new_n797), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT105), .Z(new_n947));
  NOR3_X1   g522(.A1(new_n939), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n935), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n688), .B(new_n691), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n949), .A2(new_n712), .A3(new_n715), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT103), .Z(new_n955));
  NOR2_X1   g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G8), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT120), .B1(G168), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT120), .ZN(new_n959));
  NAND3_X1  g534(.A1(G286), .A2(new_n959), .A3(G8), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n828), .A2(new_n962), .A3(new_n929), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n492), .B2(new_n496), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n964), .B2(new_n962), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2084), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n828), .A2(KEYINPUT106), .A3(new_n962), .A4(new_n929), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n933), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n969), .A2(KEYINPUT113), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n934), .B1(new_n963), .B2(new_n965), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n967), .A4(new_n968), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT96), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n492), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n488), .A2(KEYINPUT96), .A3(new_n491), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n977), .B2(new_n496), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(new_n964), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n933), .B1(new_n980), .B2(new_n931), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n734), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n961), .B1(new_n970), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT121), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n961), .B(KEYINPUT121), .C1(new_n970), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n989));
  AND2_X1   g564(.A1(new_n973), .A2(new_n982), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n969), .A2(KEYINPUT113), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n957), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n989), .B1(new_n992), .B2(new_n961), .ZN(new_n993));
  OAI21_X1  g568(.A(G8), .B1(new_n970), .B2(new_n983), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(KEYINPUT51), .A3(new_n960), .A4(new_n958), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n996), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT125), .B1(new_n996), .B2(KEYINPUT62), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n988), .A2(new_n993), .A3(new_n999), .A4(new_n995), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n828), .A2(new_n933), .A3(new_n929), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n577), .A2(new_n1004), .A3(new_n578), .A4(new_n579), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n579), .A2(new_n578), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n575), .A2(new_n576), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1008), .A2(new_n1009), .B1(new_n1010), .B2(G651), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n579), .A2(new_n578), .A3(KEYINPUT110), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1007), .B(KEYINPUT49), .C1(new_n1013), .C2(new_n1004), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1005), .B(KEYINPUT109), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1003), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT108), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1003), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(G8), .A3(new_n1001), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1019), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n966), .A2(new_n1028), .A3(new_n968), .A4(new_n933), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n828), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n980), .A2(new_n931), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n933), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n697), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n957), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT107), .B(KEYINPUT55), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G166), .A2(new_n957), .ZN(new_n1037));
  MUX2_X1   g612(.A(new_n1035), .B(new_n1036), .S(new_n1037), .Z(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n964), .B2(new_n962), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n964), .A2(new_n1040), .A3(new_n962), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n934), .B1(new_n930), .B2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1028), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n957), .B1(new_n1046), .B2(new_n1033), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1027), .B(new_n1039), .C1(new_n1038), .C2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n966), .A2(new_n968), .A3(new_n933), .ZN(new_n1049));
  INV_X1    g624(.A(G1961), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1030), .A2(new_n1031), .A3(new_n784), .A4(new_n933), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1049), .A2(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n979), .A2(new_n981), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1000), .A2(new_n1058), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n997), .A2(new_n998), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT63), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(G168), .C1(new_n970), .C2(new_n983), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1048), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT114), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1061), .C1(new_n1048), .C2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1039), .A2(KEYINPUT63), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1019), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1038), .B1(new_n1034), .B2(KEYINPUT115), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1064), .B(new_n1066), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n557), .B(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT117), .B(G1956), .Z(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n933), .B1(new_n978), .B2(new_n962), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n964), .A2(new_n1040), .A3(new_n962), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1041), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n934), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1031), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1078), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n978), .A2(new_n1090), .A3(new_n933), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1001), .A2(KEYINPUT119), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1089), .A2(new_n1049), .B1(new_n1093), .B2(new_n943), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n598), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1084), .A2(new_n1078), .A3(new_n1087), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1088), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND3_X1  g673(.A1(new_n1091), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1030), .A2(new_n1031), .A3(new_n937), .A4(new_n933), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n545), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n541), .A2(new_n544), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1103), .B(new_n1104), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1079), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n557), .B(new_n1077), .Z(new_n1109));
  AND4_X1   g684(.A1(new_n933), .A2(new_n1030), .A3(new_n1031), .A4(new_n1086), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1107), .B1(new_n1111), .B2(new_n1088), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n598), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1096), .A3(KEYINPUT61), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1106), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n598), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1097), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1052), .A2(new_n1051), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1085), .A2(KEYINPUT53), .A3(new_n784), .A4(new_n932), .ZN(new_n1124));
  AND4_X1   g699(.A1(G301), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1121), .B1(new_n1125), .B2(new_n1056), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT124), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n1121), .C1(new_n1125), .C2(new_n1056), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1053), .A2(G301), .A3(new_n1055), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1053), .A2(new_n1124), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(G171), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1048), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1120), .A2(new_n1130), .A3(new_n996), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1039), .A2(new_n1069), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1019), .A2(new_n1020), .A3(new_n704), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1007), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT111), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1002), .B1(new_n1139), .B2(KEYINPUT111), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1076), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n956), .B1(new_n1060), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n936), .A2(new_n946), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT127), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n940), .B(KEYINPUT46), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT47), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n953), .B(KEYINPUT48), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n951), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n689), .A2(new_n691), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT126), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n948), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n949), .B1(new_n1154), .B2(new_n944), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1144), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g732(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G229), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g734(.A(new_n850), .B(new_n1160), .C1(new_n925), .C2(new_n926), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


