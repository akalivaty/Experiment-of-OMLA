//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n203), .A2(new_n204), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n208), .B(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n212), .B(KEYINPUT79), .Z(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G226gat), .A2(G233gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT25), .B1(new_n219), .B2(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n225), .B2(KEYINPUT66), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n232), .A2(new_n234), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n240), .A3(new_n224), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n226), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n224), .B1(new_n219), .B2(KEYINPUT23), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT65), .B(G176gat), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n249), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n233), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n218), .B1(new_n242), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  AOI211_X1 g056(.A(new_n252), .B(new_n233), .C1(new_n248), .C2(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n221), .A2(new_n222), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT65), .B(G176gat), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n261), .B(new_n224), .C1(new_n262), .C2(new_n245), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n226), .A2(new_n239), .A3(new_n241), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n268));
  NOR2_X1   g067(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n229), .A2(new_n231), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT27), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n271), .B2(G190gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT27), .B(G183gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n259), .A2(KEYINPUT26), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n224), .B1(new_n219), .B2(new_n277), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n276), .A2(new_n278), .B1(new_n228), .B2(new_n230), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n217), .B1(new_n267), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n272), .B2(new_n274), .ZN(new_n283));
  AOI211_X1 g082(.A(KEYINPUT80), .B(new_n283), .C1(new_n256), .C2(new_n266), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n216), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n264), .B2(new_n265), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT81), .B1(new_n288), .B2(new_n215), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n264), .A2(new_n265), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n216), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n202), .B(new_n214), .C1(new_n287), .C2(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n281), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT80), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n267), .A2(new_n217), .A3(new_n281), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n286), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n301), .B2(new_n215), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT82), .B1(new_n302), .B2(new_n213), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n282), .A2(new_n284), .A3(new_n215), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n212), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n281), .B2(new_n290), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n307), .A2(KEYINPUT83), .A3(new_n216), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT83), .B1(new_n307), .B2(new_n216), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n303), .A3(new_n310), .A4(new_n314), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT30), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n295), .A2(new_n310), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n303), .A4(new_n314), .ZN(new_n321));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT0), .ZN(new_n323));
  XNOR2_X1  g122(.A(G57gat), .B(G85gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(G127gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G127gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(G113gat), .B2(G120gat), .ZN(new_n331));
  AND2_X1   g130(.A1(G113gat), .A2(G120gat), .ZN(new_n332));
  OAI22_X1  g131(.A1(new_n327), .A2(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n331), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  OR2_X1    g136(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n333), .B(KEYINPUT72), .C1(new_n336), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n340), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n335), .A4(new_n334), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(KEYINPUT85), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n355), .B2(KEYINPUT2), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(KEYINPUT2), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n346), .A3(new_n347), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(KEYINPUT84), .A3(new_n352), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n345), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(new_n364), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n341), .B2(new_n344), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT87), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n345), .A2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT86), .B(KEYINPUT3), .Z(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n364), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n375), .A2(new_n341), .A3(new_n344), .A4(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n345), .A2(new_n365), .A3(KEYINPUT4), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n374), .A2(new_n378), .A3(new_n370), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n381), .B(new_n382), .C1(new_n366), .C2(new_n368), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n371), .A2(KEYINPUT5), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(KEYINPUT89), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n325), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n382), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n370), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT39), .A3(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n325), .C1(KEYINPUT39), .C2(new_n393), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT40), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n318), .A2(new_n321), .A3(new_n391), .A4(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n212), .A2(KEYINPUT29), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n367), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n286), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n399), .B(new_n401), .C1(new_n213), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n208), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(new_n209), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n209), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n286), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n365), .B1(new_n408), .B2(new_n376), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n212), .B2(new_n402), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n404), .B1(new_n399), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  MUX2_X1   g215(.A(G22gat), .B(new_n413), .S(new_n416), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n411), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n315), .B1(new_n311), .B2(KEYINPUT37), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n311), .A2(KEYINPUT37), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n302), .A2(new_n213), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n308), .A2(new_n309), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n212), .B1(new_n425), .B2(new_n304), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT38), .B1(new_n427), .B2(KEYINPUT37), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n315), .C1(KEYINPUT37), .C2(new_n311), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n325), .B1(new_n384), .B2(new_n385), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  INV_X1    g231(.A(new_n325), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n386), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n431), .B1(new_n390), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n317), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n398), .B(new_n418), .C1(new_n423), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n341), .A2(new_n344), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n281), .B(new_n441), .C1(new_n296), .C2(new_n297), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n283), .B1(new_n256), .B2(new_n266), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n444), .A2(new_n441), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT75), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(new_n448), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g258(.A(KEYINPUT74), .B(KEYINPUT33), .C1(new_n446), .C2(new_n448), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n442), .B(new_n447), .C1(new_n443), .C2(new_n445), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT34), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n441), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n298), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n447), .A4(new_n442), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n468), .A2(KEYINPUT76), .B1(new_n449), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT76), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n463), .A2(new_n472), .A3(new_n467), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n470), .A3(new_n473), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(KEYINPUT36), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n318), .A2(new_n321), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n431), .B1(new_n434), .B2(new_n430), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n418), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n475), .B2(new_n476), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n487), .A2(new_n490), .A3(new_n435), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n438), .A2(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT13), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(G43gat), .ZN(new_n497));
  INV_X1    g296(.A(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G50gat), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(KEYINPUT93), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT15), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n504), .A2(new_n509), .A3(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n503), .B(new_n513), .C1(KEYINPUT93), .C2(new_n499), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n498), .A2(G43gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n501), .A3(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n514), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT95), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT16), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT94), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n526), .B(new_n528), .C1(new_n525), .C2(new_n524), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(KEYINPUT94), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n529), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(new_n523), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n529), .B(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n519), .A3(new_n521), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT95), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n496), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n514), .A2(new_n519), .A3(new_n542), .A4(new_n521), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n534), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n494), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n539), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n494), .A4(new_n544), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G169gat), .B(G197gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT12), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n546), .B(new_n557), .C1(new_n549), .C2(new_n550), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT104), .B(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n567), .A2(new_n572), .A3(new_n568), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n541), .A2(new_n543), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n522), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G190gat), .B(G218gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n583), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G71gat), .B(G78gat), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(G64gat), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(KEYINPUT97), .A3(G57gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n599), .B(new_n601), .C1(G57gat), .C2(new_n600), .ZN(new_n602));
  XNOR2_X1  g401(.A(G71gat), .B(G78gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n593), .A2(new_n596), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n594), .B1(new_n606), .B2(new_n591), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT101), .B(KEYINPUT19), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n532), .B1(KEYINPUT21), .B2(new_n608), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT20), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT100), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n590), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n575), .A3(new_n574), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n607), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n576), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n626), .A2(new_n628), .A3(KEYINPUT105), .A4(new_n629), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n628), .ZN(new_n642));
  INV_X1    g441(.A(new_n636), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n635), .A2(KEYINPUT106), .A3(new_n636), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n647), .A2(new_n648), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n645), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n625), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n493), .A2(new_n562), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n483), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n493), .A2(new_n562), .ZN(new_n657));
  INV_X1    g456(.A(new_n482), .ZN(new_n658));
  INV_X1    g457(.A(new_n652), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT42), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n663), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n660), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1325gat));
  AOI21_X1  g467(.A(G15gat), .B1(new_n653), .B2(new_n477), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n481), .A2(G15gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT108), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n653), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n485), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n623), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n657), .A2(new_n676), .A3(new_n589), .A4(new_n651), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n505), .A3(new_n654), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n623), .B(KEYINPUT109), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n561), .A3(new_n651), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT110), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(KEYINPUT111), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(KEYINPUT111), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n493), .B2(new_n590), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n461), .A2(new_n470), .A3(new_n473), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n473), .B1(new_n461), .B2(new_n470), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n690), .A2(new_n691), .A3(new_n478), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT36), .B1(new_n475), .B2(new_n476), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n654), .B1(new_n318), .B2(new_n321), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n418), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n317), .B(new_n431), .C1(new_n390), .C2(new_n434), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(new_n421), .B2(new_n428), .ZN(new_n698));
  INV_X1    g497(.A(new_n422), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT38), .B1(new_n699), .B2(new_n420), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n485), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n696), .B1(new_n398), .B2(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n488), .A2(KEYINPUT35), .B1(new_n491), .B2(new_n482), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n589), .B(new_n685), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n682), .B1(new_n689), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n483), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n679), .A2(new_n707), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n677), .A2(new_n509), .A3(new_n658), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n706), .B2(new_n482), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(new_n497), .B1(new_n706), .B2(new_n694), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n497), .B1(new_n475), .B2(new_n476), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n677), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n706), .B2(new_n418), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT113), .A2(KEYINPUT48), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n418), .A2(G50gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n677), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(KEYINPUT113), .A2(KEYINPUT48), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1331gat));
  NAND3_X1  g525(.A1(new_n625), .A2(new_n562), .A3(new_n650), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n493), .A2(KEYINPUT114), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT114), .B1(new_n493), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n483), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n598), .ZN(G1332gat));
  AOI21_X1  g531(.A(new_n482), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n730), .A2(KEYINPUT115), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT115), .B1(new_n730), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n730), .B2(new_n694), .ZN(new_n740));
  INV_X1    g539(.A(G71gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n477), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n418), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g546(.A1(new_n561), .A2(new_n623), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n650), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n688), .B2(new_n704), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n483), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n589), .B(new_n748), .C1(new_n702), .C2(new_n703), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n486), .A2(new_n438), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n489), .A2(new_n492), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n590), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n651), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n564), .A3(new_n654), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n752), .A2(new_n761), .ZN(G1336gat));
  AOI211_X1 g561(.A(new_n482), .B(new_n749), .C1(new_n688), .C2(new_n704), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n482), .A2(new_n651), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n565), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n755), .B2(new_n759), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n763), .A2(new_n565), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n765), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n758), .B2(new_n748), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT119), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(new_n766), .B2(new_n767), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n750), .A2(new_n658), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT118), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n776), .A2(new_n778), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(new_n763), .B2(new_n565), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n785), .A3(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n779), .A2(KEYINPUT117), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n784), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n791), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n751), .B2(new_n694), .ZN(new_n793));
  INV_X1    g592(.A(G99gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n760), .A2(new_n794), .A3(new_n477), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n760), .A2(new_n797), .A3(new_n485), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n751), .A2(new_n418), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n797), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n635), .A2(KEYINPUT106), .A3(new_n636), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT106), .B1(new_n635), .B2(new_n636), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT54), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n632), .A2(new_n643), .A3(new_n633), .A4(new_n634), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n637), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n641), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n647), .A2(new_n810), .A3(new_n648), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n635), .B2(new_n636), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n640), .B1(new_n812), .B2(new_n806), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n561), .A2(new_n809), .A3(new_n645), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n537), .A2(new_n544), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(G229gat), .A3(G233gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n537), .A2(new_n538), .A3(new_n496), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n556), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n560), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n650), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n589), .B1(new_n815), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n590), .A2(new_n824), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n814), .A2(new_n645), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n829), .A3(new_n809), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n680), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n659), .A2(new_n562), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n485), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n654), .A3(new_n482), .A4(new_n477), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n337), .A3(new_n562), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n483), .B1(new_n831), .B2(new_n832), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n487), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT121), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n658), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n561), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n835), .B1(new_n840), .B2(new_n337), .ZN(G1340gat));
  NAND4_X1  g640(.A1(new_n839), .A2(new_n338), .A3(new_n339), .A4(new_n650), .ZN(new_n842));
  OAI21_X1  g641(.A(G120gat), .B1(new_n834), .B2(new_n651), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n326), .A3(new_n623), .ZN(new_n845));
  OAI21_X1  g644(.A(G127gat), .B1(new_n834), .B2(new_n680), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  NOR2_X1   g646(.A1(new_n658), .A2(new_n590), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n328), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n834), .B2(new_n590), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n828), .A2(new_n829), .A3(new_n809), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n811), .A2(new_n813), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n559), .A2(new_n560), .B1(new_n856), .B2(new_n802), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n857), .A2(new_n829), .B1(new_n650), .B2(new_n825), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n589), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n859), .A2(new_n676), .B1(new_n562), .B2(new_n659), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n860), .B2(new_n418), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n418), .B1(new_n831), .B2(new_n832), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n658), .A2(new_n481), .A3(new_n483), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G141gat), .B1(new_n866), .B2(new_n562), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n481), .A2(new_n418), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n836), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n658), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n562), .A2(G141gat), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT58), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n676), .B1(new_n827), .B2(new_n830), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n418), .B1(new_n875), .B2(new_n832), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n865), .B1(new_n876), .B2(new_n863), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT57), .B(new_n418), .C1(new_n831), .C2(new_n832), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT122), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n864), .A3(new_n880), .A4(new_n865), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n561), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n874), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT123), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n873), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  AND2_X1   g688(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n650), .A3(new_n865), .ZN(new_n893));
  INV_X1    g692(.A(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT59), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n650), .A3(new_n881), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n894), .A2(KEYINPUT59), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(KEYINPUT124), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT124), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n870), .A2(new_n894), .A3(new_n650), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1345gat));
  NAND2_X1  g701(.A1(new_n879), .A2(new_n881), .ZN(new_n903));
  OAI21_X1  g702(.A(G155gat), .B1(new_n903), .B2(new_n680), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n870), .A2(new_n353), .A3(new_n623), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n903), .B2(new_n590), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n848), .A2(new_n354), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n869), .B2(new_n908), .ZN(G1347gat));
  AOI21_X1  g708(.A(new_n654), .B1(new_n831), .B2(new_n832), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n658), .A3(new_n487), .ZN(new_n911));
  AOI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n561), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n833), .A2(new_n483), .A3(new_n658), .A4(new_n477), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(new_n221), .A3(new_n562), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(G1348gat));
  AOI21_X1  g714(.A(G176gat), .B1(new_n911), .B2(new_n650), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n913), .A2(new_n244), .A3(new_n651), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n911), .A2(new_n273), .A3(new_n623), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT125), .Z(new_n920));
  OAI21_X1  g719(.A(new_n270), .B1(new_n913), .B2(new_n680), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n913), .B2(new_n590), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n230), .A3(new_n589), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1351gat));
  NOR3_X1   g729(.A1(new_n481), .A2(new_n654), .A3(new_n482), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n892), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(G197gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(new_n562), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n910), .A2(new_n868), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n482), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n561), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n934), .A2(new_n937), .ZN(G1352gat));
  XOR2_X1   g737(.A(KEYINPUT126), .B(G204gat), .Z(new_n939));
  NAND4_X1  g738(.A1(new_n910), .A2(new_n764), .A3(new_n868), .A4(new_n939), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT62), .Z(new_n941));
  NOR2_X1   g740(.A1(new_n932), .A2(new_n651), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n939), .ZN(G1353gat));
  INV_X1    g742(.A(new_n936), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n944), .A2(G211gat), .A3(new_n676), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n623), .B(new_n931), .C1(new_n890), .C2(new_n891), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT127), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n932), .B2(new_n590), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n590), .A2(G218gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n944), .B2(new_n952), .ZN(G1355gat));
endmodule


