

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U546 ( .A1(n531), .A2(n530), .ZN(G164) );
  AND2_X2 U547 ( .A1(n748), .A2(n576), .ZN(n615) );
  NOR2_X2 U548 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U549 ( .A(n633), .B(KEYINPUT30), .ZN(n634) );
  XNOR2_X1 U550 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U551 ( .A1(G543), .A2(G651), .ZN(n790) );
  NOR2_X1 U552 ( .A1(n524), .A2(G2105), .ZN(n891) );
  NOR2_X1 U553 ( .A1(n551), .A2(G651), .ZN(n795) );
  NAND2_X1 U554 ( .A1(G89), .A2(n790), .ZN(n510) );
  XOR2_X1 U555 ( .A(KEYINPUT4), .B(n510), .Z(n511) );
  XNOR2_X1 U556 ( .A(n511), .B(KEYINPUT73), .ZN(n513) );
  XOR2_X1 U557 ( .A(KEYINPUT0), .B(G543), .Z(n551) );
  INV_X1 U558 ( .A(G651), .ZN(n515) );
  NOR2_X1 U559 ( .A1(n551), .A2(n515), .ZN(n791) );
  NAND2_X1 U560 ( .A1(G76), .A2(n791), .ZN(n512) );
  NAND2_X1 U561 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U562 ( .A(n514), .B(KEYINPUT5), .ZN(n521) );
  NOR2_X1 U563 ( .A1(G543), .A2(n515), .ZN(n516) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n516), .Z(n794) );
  NAND2_X1 U565 ( .A1(G63), .A2(n794), .ZN(n518) );
  NAND2_X1 U566 ( .A1(G51), .A2(n795), .ZN(n517) );
  NAND2_X1 U567 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U568 ( .A(KEYINPUT6), .B(n519), .Z(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n522), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U571 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n523), .Z(n890) );
  NAND2_X1 U574 ( .A1(G138), .A2(n890), .ZN(n531) );
  INV_X1 U575 ( .A(G2104), .ZN(n524) );
  AND2_X1 U576 ( .A1(G102), .A2(n891), .ZN(n529) );
  AND2_X1 U577 ( .A1(n524), .A2(G2105), .ZN(n886) );
  NAND2_X1 U578 ( .A1(G126), .A2(n886), .ZN(n526) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U580 ( .A1(G114), .A2(n887), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U582 ( .A(KEYINPUT90), .B(n527), .ZN(n528) );
  NOR2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G64), .A2(n794), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G52), .A2(n795), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U587 ( .A(KEYINPUT65), .B(n534), .Z(n539) );
  NAND2_X1 U588 ( .A1(G90), .A2(n790), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G77), .A2(n791), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n537), .Z(n538) );
  NOR2_X1 U592 ( .A1(n539), .A2(n538), .ZN(G171) );
  NAND2_X1 U593 ( .A1(G62), .A2(n794), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G50), .A2(n795), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U596 ( .A(KEYINPUT81), .B(n542), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G88), .A2(n790), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G75), .A2(n791), .ZN(n543) );
  AND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(G303) );
  NAND2_X1 U601 ( .A1(G49), .A2(n795), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G74), .A2(G651), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT79), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n794), .A2(n550), .ZN(n553) );
  NAND2_X1 U606 ( .A1(n551), .A2(G87), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(G288) );
  XOR2_X1 U608 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n555) );
  NAND2_X1 U609 ( .A1(G73), .A2(n791), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n555), .B(n554), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G86), .A2(n790), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G61), .A2(n794), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n795), .A2(G48), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(G305) );
  NAND2_X1 U617 ( .A1(G85), .A2(n790), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G72), .A2(n791), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G60), .A2(n794), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G47), .A2(n795), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  OR2_X1 U623 ( .A1(n567), .A2(n566), .ZN(G290) );
  NAND2_X1 U624 ( .A1(G137), .A2(n890), .ZN(n569) );
  NAND2_X1 U625 ( .A1(G113), .A2(n887), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT64), .B(n570), .Z(n572) );
  NAND2_X1 U628 ( .A1(n886), .A2(G125), .ZN(n571) );
  AND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n748) );
  NOR2_X2 U630 ( .A1(G164), .A2(G1384), .ZN(n696) );
  INV_X1 U631 ( .A(n696), .ZN(n575) );
  NAND2_X1 U632 ( .A1(G101), .A2(n891), .ZN(n573) );
  XOR2_X1 U633 ( .A(KEYINPUT23), .B(n573), .Z(n747) );
  AND2_X1 U634 ( .A1(n747), .A2(G40), .ZN(n694) );
  INV_X1 U635 ( .A(n694), .ZN(n574) );
  NOR2_X1 U636 ( .A1(n615), .A2(G1961), .ZN(n577) );
  XNOR2_X1 U637 ( .A(n577), .B(KEYINPUT99), .ZN(n579) );
  XNOR2_X1 U638 ( .A(KEYINPUT25), .B(G2078), .ZN(n972) );
  NAND2_X1 U639 ( .A1(n615), .A2(n972), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n637) );
  NAND2_X1 U641 ( .A1(n637), .A2(G171), .ZN(n629) );
  NAND2_X1 U642 ( .A1(G65), .A2(n794), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G53), .A2(n795), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G91), .A2(n790), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G78), .A2(n791), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n915) );
  NAND2_X1 U649 ( .A1(n615), .A2(G2072), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT27), .ZN(n588) );
  INV_X1 U651 ( .A(n615), .ZN(n645) );
  AND2_X1 U652 ( .A1(G1956), .A2(n645), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n622) );
  NOR2_X1 U654 ( .A1(n915), .A2(n622), .ZN(n589) );
  XOR2_X1 U655 ( .A(n589), .B(KEYINPUT28), .Z(n626) );
  NAND2_X1 U656 ( .A1(G92), .A2(n790), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G79), .A2(n791), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G66), .A2(n794), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G54), .A2(n795), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n596), .Z(n926) );
  AND2_X1 U664 ( .A1(n615), .A2(G1996), .ZN(n598) );
  INV_X1 U665 ( .A(KEYINPUT26), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n598), .B(n597), .ZN(n612) );
  AND2_X1 U667 ( .A1(n645), .A2(G1341), .ZN(n610) );
  NAND2_X1 U668 ( .A1(G81), .A2(n790), .ZN(n599) );
  XOR2_X1 U669 ( .A(KEYINPUT69), .B(n599), .Z(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT12), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G68), .A2(n791), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U673 ( .A(KEYINPUT13), .B(n603), .ZN(n609) );
  NAND2_X1 U674 ( .A1(G56), .A2(n794), .ZN(n604) );
  XOR2_X1 U675 ( .A(KEYINPUT14), .B(n604), .Z(n607) );
  NAND2_X1 U676 ( .A1(n795), .A2(G43), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT70), .B(n605), .Z(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n924) );
  NOR2_X1 U680 ( .A1(n610), .A2(n924), .ZN(n611) );
  AND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U682 ( .A1(n926), .A2(n613), .ZN(n621) );
  NAND2_X1 U683 ( .A1(n613), .A2(n926), .ZN(n619) );
  INV_X1 U684 ( .A(n615), .ZN(n646) );
  NAND2_X1 U685 ( .A1(n646), .A2(G1348), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT100), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n615), .A2(G2067), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n915), .A2(n622), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U694 ( .A(KEYINPUT29), .B(n627), .Z(n628) );
  NAND2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n643) );
  INV_X1 U696 ( .A(G8), .ZN(n630) );
  NOR2_X1 U697 ( .A1(G1966), .A2(n630), .ZN(n631) );
  AND2_X1 U698 ( .A1(n645), .A2(n631), .ZN(n658) );
  NOR2_X1 U699 ( .A1(G2084), .A2(n646), .ZN(n655) );
  NOR2_X1 U700 ( .A1(n658), .A2(n655), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n632), .A2(G8), .ZN(n635) );
  INV_X1 U702 ( .A(KEYINPUT101), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n636), .A2(G168), .ZN(n639) );
  NOR2_X1 U704 ( .A1(G171), .A2(n637), .ZN(n638) );
  NOR2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n641) );
  INV_X1 U706 ( .A(KEYINPUT31), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U708 ( .A1(n643), .A2(n642), .ZN(n656) );
  NAND2_X1 U709 ( .A1(n656), .A2(G286), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n644), .B(KEYINPUT102), .ZN(n652) );
  NAND2_X1 U711 ( .A1(n645), .A2(G8), .ZN(n689) );
  NOR2_X1 U712 ( .A1(G1971), .A2(n689), .ZN(n648) );
  NOR2_X1 U713 ( .A1(G2090), .A2(n646), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U715 ( .A1(n649), .A2(G303), .ZN(n650) );
  XOR2_X1 U716 ( .A(KEYINPUT103), .B(n650), .Z(n651) );
  NAND2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U718 ( .A1(n653), .A2(G8), .ZN(n654) );
  XNOR2_X1 U719 ( .A(n654), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U720 ( .A1(G8), .A2(n655), .ZN(n660) );
  INV_X1 U721 ( .A(n656), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n680) );
  NAND2_X1 U724 ( .A1(G288), .A2(G1976), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT105), .B(n661), .Z(n920) );
  AND2_X1 U726 ( .A1(n680), .A2(n920), .ZN(n663) );
  INV_X1 U727 ( .A(KEYINPUT33), .ZN(n662) );
  AND2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n679), .A2(n664), .ZN(n670) );
  INV_X1 U730 ( .A(n920), .ZN(n667) );
  NOR2_X1 U731 ( .A1(G1976), .A2(G288), .ZN(n912) );
  NOR2_X1 U732 ( .A1(G1971), .A2(G303), .ZN(n911) );
  XNOR2_X1 U733 ( .A(KEYINPUT104), .B(n911), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n912), .A2(n665), .ZN(n666) );
  OR2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  OR2_X1 U736 ( .A1(KEYINPUT33), .A2(n668), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  INV_X1 U738 ( .A(n689), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n671), .A2(n672), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n912), .A2(n672), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n673), .A2(KEYINPUT33), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(KEYINPUT106), .ZN(n678) );
  XNOR2_X1 U744 ( .A(KEYINPUT107), .B(G1981), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(G305), .ZN(n929) );
  NAND2_X1 U746 ( .A1(n678), .A2(n929), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n683) );
  NOR2_X1 U748 ( .A1(G2090), .A2(G303), .ZN(n681) );
  NAND2_X1 U749 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n689), .A2(n684), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n693) );
  NOR2_X1 U753 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n687), .B(KEYINPUT24), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n688), .B(KEYINPUT97), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n691), .B(KEYINPUT98), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n718) );
  NAND2_X1 U759 ( .A1(n748), .A2(n694), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n743) );
  NAND2_X1 U761 ( .A1(G95), .A2(n891), .ZN(n703) );
  NAND2_X1 U762 ( .A1(G119), .A2(n886), .ZN(n698) );
  NAND2_X1 U763 ( .A1(G107), .A2(n887), .ZN(n697) );
  NAND2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U765 ( .A1(G131), .A2(n890), .ZN(n699) );
  XNOR2_X1 U766 ( .A(KEYINPUT93), .B(n699), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT94), .ZN(n866) );
  NAND2_X1 U770 ( .A1(n866), .A2(G1991), .ZN(n715) );
  NAND2_X1 U771 ( .A1(G129), .A2(n886), .ZN(n706) );
  NAND2_X1 U772 ( .A1(G117), .A2(n887), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n707), .B(KEYINPUT95), .ZN(n709) );
  NAND2_X1 U775 ( .A1(G141), .A2(n890), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n891), .A2(G105), .ZN(n710) );
  XOR2_X1 U778 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U780 ( .A(KEYINPUT96), .B(n713), .Z(n869) );
  NAND2_X1 U781 ( .A1(n869), .A2(G1996), .ZN(n714) );
  NAND2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n1003) );
  NAND2_X1 U783 ( .A1(n743), .A2(n1003), .ZN(n732) );
  XNOR2_X1 U784 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U785 ( .A1(n743), .A2(n919), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n732), .A2(n716), .ZN(n717) );
  NOR2_X2 U787 ( .A1(n718), .A2(n717), .ZN(n730) );
  NAND2_X1 U788 ( .A1(G128), .A2(n886), .ZN(n720) );
  NAND2_X1 U789 ( .A1(G116), .A2(n887), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U791 ( .A(n721), .B(KEYINPUT35), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n890), .A2(G140), .ZN(n722) );
  XOR2_X1 U793 ( .A(KEYINPUT91), .B(n722), .Z(n724) );
  NAND2_X1 U794 ( .A1(n891), .A2(G104), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U796 ( .A(KEYINPUT34), .B(n725), .Z(n726) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U798 ( .A(n728), .B(KEYINPUT36), .Z(n867) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n740) );
  OR2_X1 U800 ( .A1(n867), .A2(n740), .ZN(n729) );
  XOR2_X1 U801 ( .A(KEYINPUT92), .B(n729), .Z(n1007) );
  NAND2_X1 U802 ( .A1(n743), .A2(n1007), .ZN(n738) );
  NAND2_X1 U803 ( .A1(n730), .A2(n738), .ZN(n731) );
  XNOR2_X1 U804 ( .A(n731), .B(KEYINPUT108), .ZN(n745) );
  NOR2_X1 U805 ( .A1(G1996), .A2(n869), .ZN(n996) );
  INV_X1 U806 ( .A(n732), .ZN(n735) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n866), .ZN(n994) );
  NOR2_X1 U809 ( .A1(n733), .A2(n994), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n996), .A2(n736), .ZN(n737) );
  XNOR2_X1 U812 ( .A(KEYINPUT39), .B(n737), .ZN(n739) );
  NAND2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n867), .A2(n740), .ZN(n1008) );
  NAND2_X1 U815 ( .A1(n741), .A2(n1008), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U818 ( .A(n746), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U819 ( .A1(n748), .A2(n747), .ZN(G160) );
  XOR2_X1 U820 ( .A(G2430), .B(G2451), .Z(n750) );
  XNOR2_X1 U821 ( .A(KEYINPUT109), .B(G2443), .ZN(n749) );
  XNOR2_X1 U822 ( .A(n750), .B(n749), .ZN(n757) );
  XOR2_X1 U823 ( .A(G2435), .B(G2446), .Z(n752) );
  XNOR2_X1 U824 ( .A(G2427), .B(G2454), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U826 ( .A(n753), .B(G2438), .Z(n755) );
  XNOR2_X1 U827 ( .A(G1341), .B(G1348), .ZN(n754) );
  XNOR2_X1 U828 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n757), .B(n756), .ZN(n758) );
  AND2_X1 U830 ( .A1(n758), .A2(G14), .ZN(G401) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(G82), .ZN(G220) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n761) );
  XNOR2_X1 U837 ( .A(G223), .B(KEYINPUT67), .ZN(n833) );
  NAND2_X1 U838 ( .A1(G567), .A2(n833), .ZN(n760) );
  XNOR2_X1 U839 ( .A(n761), .B(n760), .ZN(G234) );
  INV_X1 U840 ( .A(G860), .ZN(n770) );
  OR2_X1 U841 ( .A1(n924), .A2(n770), .ZN(n762) );
  XOR2_X1 U842 ( .A(KEYINPUT71), .B(n762), .Z(G153) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  NAND2_X1 U844 ( .A1(G301), .A2(G868), .ZN(n763) );
  XNOR2_X1 U845 ( .A(n763), .B(KEYINPUT72), .ZN(n765) );
  INV_X1 U846 ( .A(G868), .ZN(n812) );
  INV_X1 U847 ( .A(n926), .ZN(n774) );
  NAND2_X1 U848 ( .A1(n812), .A2(n774), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(G284) );
  INV_X1 U850 ( .A(n915), .ZN(G299) );
  XNOR2_X1 U851 ( .A(KEYINPUT74), .B(n812), .ZN(n766) );
  NOR2_X1 U852 ( .A1(G286), .A2(n766), .ZN(n767) );
  XOR2_X1 U853 ( .A(KEYINPUT75), .B(n767), .Z(n769) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n770), .A2(G559), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n771), .A2(n926), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT76), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT16), .B(n773), .ZN(G148) );
  NOR2_X1 U860 ( .A1(n774), .A2(n812), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT77), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G559), .A2(n776), .ZN(n778) );
  NOR2_X1 U863 ( .A1(G868), .A2(n924), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U865 ( .A1(n886), .A2(G123), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G135), .A2(n890), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(KEYINPUT78), .B(n782), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G111), .A2(n887), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G99), .A2(n891), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n993) );
  XNOR2_X1 U874 ( .A(n993), .B(G2096), .ZN(n788) );
  INV_X1 U875 ( .A(G2100), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U877 ( .A1(n926), .A2(G559), .ZN(n809) );
  XNOR2_X1 U878 ( .A(n924), .B(n809), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n789), .A2(G860), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G67), .A2(n794), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G55), .A2(n795), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n811) );
  XOR2_X1 U887 ( .A(n800), .B(n811), .Z(G145) );
  XOR2_X1 U888 ( .A(G290), .B(n924), .Z(n801) );
  XOR2_X1 U889 ( .A(n811), .B(n801), .Z(n806) );
  XOR2_X1 U890 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n803) );
  XNOR2_X1 U891 ( .A(n915), .B(KEYINPUT83), .ZN(n802) );
  XNOR2_X1 U892 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U893 ( .A(G305), .B(n804), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(G288), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n808), .B(G303), .ZN(n901) );
  XNOR2_X1 U897 ( .A(n809), .B(n901), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n810), .A2(G868), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U906 ( .A1(G2072), .A2(n819), .ZN(G158) );
  XOR2_X1 U907 ( .A(KEYINPUT85), .B(G44), .Z(n820) );
  XNOR2_X1 U908 ( .A(KEYINPUT3), .B(n820), .ZN(G218) );
  XOR2_X1 U909 ( .A(KEYINPUT66), .B(G132), .Z(G219) );
  NAND2_X1 U910 ( .A1(G120), .A2(G69), .ZN(n821) );
  NOR2_X1 U911 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n822), .A2(G108), .ZN(n823) );
  XNOR2_X1 U913 ( .A(n823), .B(KEYINPUT88), .ZN(n839) );
  NAND2_X1 U914 ( .A1(G567), .A2(n839), .ZN(n830) );
  NOR2_X1 U915 ( .A1(G219), .A2(G220), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT86), .B(n824), .Z(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT22), .ZN(n826) );
  NOR2_X1 U918 ( .A1(G218), .A2(n826), .ZN(n827) );
  XOR2_X1 U919 ( .A(KEYINPUT87), .B(n827), .Z(n828) );
  NAND2_X1 U920 ( .A1(G96), .A2(n828), .ZN(n838) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n838), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n857) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n831) );
  XOR2_X1 U924 ( .A(KEYINPUT89), .B(n831), .Z(n832) );
  NOR2_X1 U925 ( .A1(n857), .A2(n832), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n837), .A2(G36), .ZN(G176) );
  INV_X1 U927 ( .A(G303), .ZN(G166) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  XOR2_X1 U930 ( .A(KEYINPUT110), .B(n834), .Z(n835) );
  NAND2_X1 U931 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U934 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1956), .B(G1961), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U952 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1976), .B(G1971), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1981), .Z(n854) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U959 ( .A(KEYINPUT112), .B(n857), .Z(G319) );
  NAND2_X1 U960 ( .A1(G124), .A2(n886), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G112), .A2(n887), .ZN(n859) );
  XOR2_X1 U963 ( .A(KEYINPUT113), .B(n859), .Z(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G136), .A2(n890), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G100), .A2(n891), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U968 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U969 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(n993), .ZN(n880) );
  XNOR2_X1 U971 ( .A(G164), .B(n869), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G139), .A2(n890), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G103), .A2(n891), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT115), .B(n872), .Z(n877) );
  NAND2_X1 U976 ( .A1(G127), .A2(n886), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G115), .A2(n887), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n989) );
  XNOR2_X1 U981 ( .A(n878), .B(n989), .ZN(n879) );
  XOR2_X1 U982 ( .A(n880), .B(n879), .Z(n885) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U984 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U985 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U986 ( .A(G162), .B(n883), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n899) );
  NAND2_X1 U988 ( .A1(G130), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G118), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U999 ( .A(n901), .B(G286), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G171), .B(n926), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT49), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n906), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n907), .A2(G319), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT117), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1012 ( .A(G171), .B(G1961), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n923) );
  XNOR2_X1 U1015 ( .A(n915), .B(G1956), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n936) );
  XNOR2_X1 U1021 ( .A(G1341), .B(KEYINPUT123), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(n926), .B(G1348), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n934) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G168), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT57), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT122), .B(n932), .Z(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(n937), .B(KEYINPUT124), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G16), .B(KEYINPUT121), .Z(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT56), .B(n938), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n1017) );
  XNOR2_X1 U1035 ( .A(G21), .B(G1966), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(KEYINPUT127), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(G20), .B(G1956), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n942), .B(KEYINPUT125), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .Z(n943) );
  XNOR2_X1 U1040 ( .A(G4), .B(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G19), .B(G1341), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT126), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1047 ( .A(KEYINPUT60), .B(n951), .Z(n953) );
  XNOR2_X1 U1048 ( .A(G1961), .B(G5), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G1976), .B(G23), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n959) );
  XOR2_X1 U1054 ( .A(G1986), .B(G24), .Z(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT61), .B(n963), .ZN(n965) );
  INV_X1 U1059 ( .A(G16), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(G11), .ZN(n1015) );
  XOR2_X1 U1062 ( .A(KEYINPUT119), .B(G34), .Z(n968) );
  XNOR2_X1 U1063 ( .A(G2084), .B(KEYINPUT54), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(n968), .B(n967), .ZN(n985) );
  XOR2_X1 U1065 ( .A(G2090), .B(G35), .Z(n983) );
  XOR2_X1 U1066 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1067 ( .A1(n969), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G26), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(G33), .B(G2072), .ZN(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n977) );
  XOR2_X1 U1071 ( .A(n972), .B(G27), .Z(n975) );
  INV_X1 U1072 ( .A(G1996), .ZN(n973) );
  XOR2_X1 U1073 ( .A(n973), .B(G32), .Z(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1077 ( .A(KEYINPUT118), .B(n980), .Z(n981) );
  XNOR2_X1 U1078 ( .A(n981), .B(KEYINPUT53), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(KEYINPUT120), .B(n986), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(G29), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(n988), .B(KEYINPUT55), .ZN(n1013) );
  XOR2_X1 U1084 ( .A(G2072), .B(n989), .Z(n991) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT50), .B(n992), .ZN(n1005) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G160), .B(G2084), .Z(n999) );
  XOR2_X1 U1090 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(KEYINPUT51), .B(n997), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(G29), .A2(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

