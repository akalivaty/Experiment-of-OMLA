//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n208), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(KEYINPUT26), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n210), .B(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(KEYINPUT26), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n219));
  OAI221_X1 g018(.A(new_n209), .B1(KEYINPUT28), .B2(new_n208), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n225), .A2(new_n207), .A3(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(KEYINPUT24), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g027(.A(new_n222), .B1(new_n221), .B2(new_n217), .C1(new_n224), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n223), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT25), .B1(new_n210), .B2(KEYINPUT23), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n220), .B(new_n230), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G113gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT67), .B(G120gat), .Z(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  AOI211_X1 g040(.A(KEYINPUT1), .B(new_n236), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n241), .B2(new_n240), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n236), .B1(KEYINPUT1), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n234), .B(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(G227gat), .A3(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n205), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n247), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT34), .ZN(new_n252));
  NAND2_X1  g051(.A1(G227gat), .A2(G233gat), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n250), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(KEYINPUT32), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n258), .B1(new_n262), .B2(new_n256), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n202), .B1(new_n264), .B2(KEYINPUT70), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT36), .ZN(new_n268));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(KEYINPUT22), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n270), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G155gat), .B(G162gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(G155gat), .B2(G162gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n279), .B(new_n278), .C1(new_n283), .C2(new_n282), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n277), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n286), .A2(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(new_n275), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n295), .A2(new_n269), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n291), .B1(new_n295), .B2(new_n269), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n293), .A2(new_n299), .B1(G228gat), .B2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n292), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G228gat), .ZN(new_n303));
  INV_X1    g102(.A(G233gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n289), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT77), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n300), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G22gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT31), .B(G50gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n300), .ZN(new_n320));
  INV_X1    g119(.A(new_n310), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n309), .B1(new_n302), .B2(new_n306), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n312), .B1(new_n323), .B2(KEYINPUT78), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n324), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n319), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(G22gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n317), .B1(new_n331), .B2(new_n313), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335));
  AND2_X1   g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n234), .B2(new_n291), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n336), .B2(new_n234), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(new_n277), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n335), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n339), .A2(new_n343), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n246), .B(new_n294), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n246), .A2(new_n294), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT4), .B1(new_n246), .B2(new_n294), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n349), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n246), .A2(new_n290), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT73), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n351), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT74), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n359), .B(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n349), .A3(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n366), .B2(new_n351), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n369), .A3(new_n353), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n355), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n365), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI22_X1  g173(.A1(new_n362), .A2(new_n367), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OAI221_X1 g181(.A(new_n379), .B1(new_n372), .B2(new_n374), .C1(new_n362), .C2(new_n367), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n346), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n265), .B(new_n268), .C1(new_n334), .C2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n374), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n361), .A2(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n363), .A3(new_n351), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n382), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n375), .A2(new_n380), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT80), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n342), .B1(new_n339), .B2(KEYINPUT37), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(KEYINPUT37), .B2(new_n339), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT38), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n345), .B1(new_n399), .B2(KEYINPUT38), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n395), .A2(new_n397), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n324), .A2(new_n327), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT79), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n318), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n332), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT40), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n372), .A2(new_n350), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n348), .A2(new_n350), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n410), .A2(KEYINPUT39), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n379), .B1(new_n410), .B2(KEYINPUT39), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n346), .A2(new_n381), .A3(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n412), .A2(new_n413), .A3(new_n409), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n387), .B1(new_n403), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n391), .A2(new_n382), .A3(new_n379), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT6), .B1(new_n375), .B2(new_n380), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n383), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n397), .B1(new_n422), .B2(new_n396), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n266), .B1(new_n330), .B2(new_n333), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  INV_X1    g224(.A(new_n346), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n334), .A2(new_n394), .A3(new_n426), .A4(new_n264), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n427), .A2(new_n428), .B1(KEYINPUT35), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n346), .B(new_n266), .C1(new_n330), .C2(new_n333), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n431), .A2(KEYINPUT81), .A3(new_n425), .A4(new_n423), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n419), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G113gat), .B(G141gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(G197gat), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT11), .B(G169gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n437), .B(KEYINPUT12), .Z(new_n438));
  NAND2_X1  g237(.A1(G229gat), .A2(G233gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT13), .Z(new_n440));
  NOR2_X1   g239(.A1(G43gat), .A2(G50gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g242(.A1(G43gat), .A2(G50gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT14), .ZN(new_n446));
  INV_X1    g245(.A(G29gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n449));
  AOI21_X1  g248(.A(G36gat), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n444), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  INV_X1    g254(.A(new_n444), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n441), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n457), .A3(KEYINPUT15), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G36gat), .ZN(new_n460));
  AND2_X1   g259(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n451), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT15), .A3(new_n454), .A4(new_n457), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468));
  INV_X1    g267(.A(G8gat), .ZN(new_n469));
  INV_X1    g268(.A(G15gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G22gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n312), .A2(G15gat), .ZN(new_n472));
  INV_X1    g271(.A(G1gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(G1gat), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n468), .B(new_n469), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g280(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(new_n475), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT87), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n483), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n467), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT87), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT87), .B1(new_n478), .B2(new_n483), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n489), .A2(new_n490), .A3(new_n466), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n440), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT89), .B(new_n440), .C1(new_n488), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI211_X1 g295(.A(KEYINPUT84), .B(KEYINPUT17), .C1(new_n459), .C2(new_n465), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n459), .A2(new_n465), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT86), .B(new_n485), .C1(new_n497), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n491), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n466), .A2(new_n499), .A3(new_n500), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n502), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT86), .B1(new_n508), .B2(new_n485), .ZN(new_n509));
  INV_X1    g308(.A(new_n439), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n496), .B1(new_n511), .B2(KEYINPUT18), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n504), .A2(new_n505), .ZN(new_n513));
  INV_X1    g312(.A(new_n509), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(KEYINPUT18), .A3(new_n514), .A4(new_n439), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT18), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n438), .B1(new_n519), .B2(KEYINPUT82), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(new_n512), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT82), .ZN(new_n524));
  INV_X1    g323(.A(new_n438), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n433), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n533), .B(new_n532), .C1(new_n530), .C2(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT92), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(KEYINPUT91), .A2(G85gat), .ZN(new_n545));
  INV_X1    g344(.A(G92gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(KEYINPUT91), .A2(G85gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(KEYINPUT92), .A3(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(KEYINPUT8), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(KEYINPUT90), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n544), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n558), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n561), .A2(new_n562), .A3(new_n543), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n540), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n551), .A2(new_n559), .A3(new_n544), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n543), .B1(new_n561), .B2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n539), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n565), .A4(new_n568), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n565), .B(new_n539), .C1(new_n566), .C2(new_n567), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n564), .A2(new_n568), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G120gat), .B(G148gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT95), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n577), .A2(new_n580), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n579), .B1(new_n590), .B2(new_n572), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n579), .B2(new_n578), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n539), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G127gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n487), .A2(new_n484), .B1(KEYINPUT21), .B2(new_n540), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n602), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n566), .A2(new_n567), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n467), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n507), .B2(new_n502), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n610), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n529), .A2(new_n595), .A3(new_n607), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n422), .A2(KEYINPUT97), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n422), .A2(KEYINPUT97), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT98), .B(G1gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1324gat));
  XOR2_X1   g433(.A(KEYINPUT16), .B(G8gat), .Z(new_n635));
  OAI211_X1 g434(.A(new_n346), .B(new_n635), .C1(new_n626), .C2(new_n627), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(G8gat), .B1(new_n628), .B2(new_n426), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n639), .A2(new_n636), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n640), .B2(new_n637), .ZN(G1325gat));
  AOI21_X1  g440(.A(new_n628), .B1(new_n265), .B2(new_n268), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n264), .A2(new_n470), .ZN(new_n643));
  OAI22_X1  g442(.A1(new_n642), .A2(new_n470), .B1(new_n628), .B2(new_n643), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n334), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(new_n607), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n595), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n623), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n529), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n631), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n447), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT45), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n433), .B2(new_n623), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n396), .B1(new_n384), .B2(new_n385), .ZN(new_n658));
  INV_X1    g457(.A(new_n397), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n425), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n426), .B(new_n264), .C1(new_n407), .C2(new_n332), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n428), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n429), .A2(KEYINPUT35), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n432), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n418), .A2(new_n403), .ZN(new_n665));
  INV_X1    g464(.A(new_n387), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n623), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n528), .A2(new_n649), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n631), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n673), .ZN(G1328gat));
  NOR3_X1   g473(.A1(new_n651), .A2(G36gat), .A3(new_n426), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT99), .B(KEYINPUT46), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n672), .B2(new_n426), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(G43gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n652), .A2(new_n680), .A3(new_n264), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n265), .A2(new_n268), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n657), .A2(new_n682), .A3(new_n669), .A4(new_n671), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT101), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n681), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT47), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n689), .B(new_n691), .ZN(G1330gat));
  NOR3_X1   g491(.A1(new_n651), .A2(G50gat), .A3(new_n334), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n670), .A2(new_n408), .A3(new_n671), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G50gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n664), .A2(new_n667), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n527), .A2(new_n648), .A3(new_n622), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n594), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n631), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n426), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  AND2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(G1333gat));
  XNOR2_X1  g510(.A(new_n264), .B(KEYINPUT104), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n682), .A2(G71gat), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n713), .A2(G71gat), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g515(.A1(new_n704), .A2(new_n334), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT105), .B(G78gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n527), .A2(new_n607), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n668), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT106), .B1(new_n433), .B2(new_n623), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n545), .A2(new_n547), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n631), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n727), .A2(new_n728), .A3(new_n594), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n720), .A2(new_n594), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n670), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n729), .B1(new_n734), .B2(new_n631), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT107), .ZN(G1336gat));
  AND2_X1   g536(.A1(new_n727), .A2(new_n728), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n426), .A2(G92gat), .A3(new_n595), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n734), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n546), .B1(new_n741), .B2(new_n346), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT52), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT108), .B1(new_n746), .B2(KEYINPUT51), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n723), .B2(new_n724), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n723), .A2(new_n724), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n746), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n748), .B1(new_n751), .B2(new_n726), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n745), .B1(new_n752), .B2(new_n739), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n750), .B2(new_n746), .ZN(new_n754));
  INV_X1    g553(.A(new_n739), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n754), .A2(KEYINPUT110), .A3(new_n748), .A4(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n753), .A2(new_n756), .A3(new_n742), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n744), .B1(new_n757), .B2(new_n758), .ZN(G1337gat));
  INV_X1    g558(.A(G99gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n682), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n738), .A2(new_n760), .A3(new_n264), .A4(new_n594), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1338gat));
  NOR3_X1   g565(.A1(new_n334), .A2(G106gat), .A3(new_n595), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n727), .A2(new_n728), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n670), .A2(new_n408), .A3(new_n733), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT112), .ZN(new_n771));
  OAI21_X1  g570(.A(G106gat), .B1(new_n770), .B2(KEYINPUT112), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n768), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n752), .A2(new_n767), .B1(G106gat), .B2(new_n770), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n769), .B2(new_n774), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n701), .A2(new_n595), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n590), .A2(new_n579), .A3(new_n572), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n577), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n779));
  AOI21_X1  g578(.A(new_n584), .B1(new_n591), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT55), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n589), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n783), .A2(KEYINPUT115), .A3(new_n589), .A4(new_n784), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n778), .A2(new_n780), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n789), .A2(KEYINPUT55), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n785), .B2(new_n786), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT116), .A3(new_n788), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n527), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n519), .A2(new_n525), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n439), .B1(new_n513), .B2(new_n514), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n488), .A2(new_n491), .A3(new_n440), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n437), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n594), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n798), .A2(new_n622), .A3(new_n801), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n804), .A3(new_n796), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n793), .A2(KEYINPUT117), .A3(new_n804), .A4(new_n796), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n623), .A2(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n776), .B1(new_n809), .B2(new_n607), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n653), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n431), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n527), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G113gat), .ZN(G1340gat));
  NOR2_X1   g615(.A1(new_n813), .A2(new_n595), .ZN(new_n817));
  MUX2_X1   g616(.A(G120gat), .B(new_n239), .S(new_n817), .Z(G1341gat));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n607), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n346), .A2(new_n623), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT118), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n812), .A2(new_n424), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT119), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n813), .B2(new_n623), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n826), .B(new_n827), .C1(KEYINPUT56), .C2(new_n824), .ZN(G1343gat));
  OR2_X1    g627(.A1(new_n631), .A2(new_n682), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n346), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n520), .A2(new_n526), .A3(new_n790), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n831), .B(new_n802), .C1(new_n832), .C2(new_n785), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n623), .ZN(new_n834));
  INV_X1    g633(.A(new_n785), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n520), .A3(new_n526), .A4(new_n790), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n831), .B1(new_n836), .B2(new_n802), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AND4_X1   g638(.A1(KEYINPUT116), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n795), .B2(new_n788), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n842), .B2(new_n804), .ZN(new_n843));
  INV_X1    g642(.A(new_n808), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(KEYINPUT122), .A3(new_n648), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n838), .B1(new_n807), .B2(new_n808), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n607), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n776), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n334), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n810), .B2(new_n408), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(KEYINPUT120), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n856), .B(KEYINPUT57), .C1(new_n810), .C2(new_n408), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n830), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n527), .A2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n810), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n334), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n830), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n528), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n858), .A2(new_n859), .B1(new_n863), .B2(G141gat), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n795), .A2(new_n804), .A3(new_n788), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n607), .B1(new_n839), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n868), .B1(new_n595), .B2(new_n701), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n851), .B1(new_n869), .B2(new_n334), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n810), .A2(KEYINPUT57), .A3(new_n408), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n594), .A3(new_n830), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n866), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n594), .B(new_n830), .C1(new_n855), .C2(new_n857), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n866), .A2(G148gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT123), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n874), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n862), .A2(G148gat), .A3(new_n595), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT124), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884));
  INV_X1    g683(.A(new_n882), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n875), .A2(new_n879), .A3(new_n876), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n884), .B(new_n885), .C1(new_n888), .C2(new_n874), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(G1345gat));
  OAI21_X1  g689(.A(G155gat), .B1(new_n858), .B2(new_n648), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n648), .A2(G155gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n862), .B2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n858), .B2(new_n623), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n829), .A2(G162gat), .A3(new_n822), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n861), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n860), .A2(new_n653), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n424), .A2(new_n346), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT125), .Z(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n527), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n631), .A2(new_n346), .ZN(new_n904));
  OR4_X1    g703(.A1(new_n408), .A2(new_n860), .A3(new_n712), .A4(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n528), .A2(new_n212), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n213), .A3(new_n594), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n594), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n213), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n905), .B2(new_n648), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n902), .A2(new_n206), .A3(new_n607), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n902), .A2(new_n207), .A3(new_n622), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n906), .A2(new_n622), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n919));
  AND4_X1   g718(.A1(KEYINPUT126), .A2(new_n918), .A3(new_n919), .A4(G190gat), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n207), .B1(new_n921), .B2(KEYINPUT61), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n918), .A2(new_n922), .B1(KEYINPUT126), .B2(new_n919), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n917), .B1(new_n920), .B2(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n682), .A2(new_n334), .A3(new_n426), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n898), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n527), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n682), .B(new_n904), .C1(new_n870), .C2(new_n871), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n527), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n926), .A2(G204gat), .A3(new_n595), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n929), .A2(new_n594), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1353gat));
  AOI21_X1  g735(.A(new_n272), .B1(new_n929), .B2(new_n607), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT63), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n272), .A3(new_n607), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1354gat));
  OAI21_X1  g739(.A(new_n273), .B1(new_n926), .B2(new_n623), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT127), .Z(new_n942));
  NOR2_X1   g741(.A1(new_n623), .A2(new_n273), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n929), .B2(new_n943), .ZN(G1355gat));
endmodule


