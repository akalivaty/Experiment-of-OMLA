

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801;

  NOR2_X1 U383 ( .A1(n616), .A2(n634), .ZN(n619) );
  NAND2_X1 U384 ( .A1(n649), .A2(n570), .ZN(n586) );
  XNOR2_X1 U385 ( .A(n410), .B(n574), .ZN(n591) );
  INV_X1 U386 ( .A(n744), .ZN(n401) );
  NOR2_X1 U387 ( .A1(n667), .A2(n741), .ZN(n744) );
  AND2_X2 U388 ( .A1(n405), .A2(n404), .ZN(n394) );
  NOR2_X2 U389 ( .A1(n627), .A2(n612), .ZN(n611) );
  NOR2_X2 U390 ( .A1(n801), .A2(n799), .ZN(n622) );
  XNOR2_X2 U391 ( .A(n528), .B(n529), .ZN(n683) );
  XNOR2_X2 U392 ( .A(n520), .B(G134), .ZN(n528) );
  OR2_X2 U393 ( .A1(n793), .A2(n381), .ZN(n440) );
  NAND2_X1 U394 ( .A1(n539), .A2(n377), .ZN(n565) );
  NAND2_X1 U395 ( .A1(n583), .A2(n582), .ZN(n420) );
  NAND2_X1 U396 ( .A1(n569), .A2(n761), .ZN(n766) );
  NOR2_X1 U397 ( .A1(n364), .A2(n466), .ZN(n798) );
  AND2_X1 U398 ( .A1(n390), .A2(n795), .ZN(n364) );
  BUF_X1 U399 ( .A(n591), .Z(n365) );
  XNOR2_X1 U400 ( .A(n465), .B(n464), .ZN(n801) );
  NAND2_X1 U401 ( .A1(n411), .A2(n625), .ZN(n410) );
  NOR2_X1 U402 ( .A1(n718), .A2(n373), .ZN(n590) );
  XNOR2_X1 U403 ( .A(n562), .B(n561), .ZN(n681) );
  NAND2_X1 U404 ( .A1(n571), .A2(n527), .ZN(n451) );
  NOR2_X1 U405 ( .A1(n604), .A2(n614), .ZN(n605) );
  INV_X1 U406 ( .A(n749), .ZN(n612) );
  XNOR2_X1 U407 ( .A(n624), .B(KEYINPUT38), .ZN(n749) );
  OR2_X1 U408 ( .A1(n441), .A2(n438), .ZN(n376) );
  XNOR2_X1 U409 ( .A(n764), .B(KEYINPUT6), .ZN(n635) );
  XNOR2_X1 U410 ( .A(n538), .B(G472), .ZN(n764) );
  XNOR2_X1 U411 ( .A(n545), .B(n546), .ZN(n712) );
  NOR2_X1 U412 ( .A1(n651), .A2(n379), .ZN(n439) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(n661), .Z(n662) );
  XNOR2_X1 U414 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n574) );
  NOR2_X1 U415 ( .A1(G902), .A2(G237), .ZN(n487) );
  INV_X1 U416 ( .A(KEYINPUT64), .ZN(n480) );
  NAND2_X1 U417 ( .A1(n394), .A2(n402), .ZN(n360) );
  NAND2_X1 U418 ( .A1(n394), .A2(n402), .ZN(n666) );
  NAND2_X1 U419 ( .A1(n539), .A2(n361), .ZN(n562) );
  AND2_X1 U420 ( .A1(n635), .A2(n560), .ZN(n361) );
  NAND2_X1 U421 ( .A1(n793), .A2(n371), .ZN(n362) );
  XNOR2_X1 U422 ( .A(G122), .B(G104), .ZN(n363) );
  NAND2_X1 U423 ( .A1(n793), .A2(n371), .ZN(n441) );
  XNOR2_X1 U424 ( .A(G122), .B(G104), .ZN(n503) );
  NAND2_X1 U425 ( .A1(n576), .A2(n575), .ZN(n407) );
  NAND2_X1 U426 ( .A1(n539), .A2(n635), .ZN(n366) );
  XNOR2_X2 U427 ( .A(n479), .B(n531), .ZN(n698) );
  XNOR2_X1 U428 ( .A(n367), .B(n368), .ZN(n673) );
  NOR2_X1 U429 ( .A1(n668), .A2(n399), .ZN(n367) );
  XOR2_X1 U430 ( .A(n670), .B(n669), .Z(n368) );
  AND2_X1 U431 ( .A1(n595), .A2(n452), .ZN(n403) );
  XNOR2_X2 U432 ( .A(n637), .B(KEYINPUT19), .ZN(n629) );
  NAND2_X2 U433 ( .A1(n426), .A2(n425), .ZN(n637) );
  NOR2_X2 U434 ( .A1(n629), .A2(n499), .ZN(n501) );
  XNOR2_X2 U435 ( .A(n698), .B(n486), .ZN(n793) );
  NAND2_X1 U436 ( .A1(n450), .A2(n413), .ZN(n412) );
  NOR2_X1 U437 ( .A1(n582), .A2(n573), .ZN(n625) );
  XNOR2_X1 U438 ( .A(n422), .B(G478), .ZN(n583) );
  NAND2_X1 U439 ( .A1(n423), .A2(n554), .ZN(n422) );
  XNOR2_X1 U440 ( .A(n417), .B(n433), .ZN(n644) );
  INV_X1 U441 ( .A(KEYINPUT77), .ZN(n433) );
  INV_X1 U442 ( .A(n721), .ZN(n436) );
  INV_X1 U443 ( .A(n739), .ZN(n656) );
  XNOR2_X1 U444 ( .A(n392), .B(n559), .ZN(n569) );
  XNOR2_X1 U445 ( .A(n558), .B(n557), .ZN(n559) );
  NOR2_X1 U446 ( .A1(G953), .A2(G237), .ZN(n530) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n508) );
  XNOR2_X1 U448 ( .A(G131), .B(G143), .ZN(n504) );
  XOR2_X1 U449 ( .A(G140), .B(G113), .Z(n502) );
  INV_X1 U450 ( .A(n586), .ZN(n459) );
  NOR2_X1 U451 ( .A1(n635), .A2(n461), .ZN(n445) );
  NOR2_X1 U452 ( .A1(n389), .A2(n379), .ZN(n388) );
  NAND2_X1 U453 ( .A1(n454), .A2(n403), .ZN(n402) );
  NAND2_X1 U454 ( .A1(n407), .A2(n577), .ZN(n454) );
  XNOR2_X1 U455 ( .A(n544), .B(n543), .ZN(n546) );
  INV_X1 U456 ( .A(KEYINPUT81), .ZN(n432) );
  AND2_X1 U457 ( .A1(n458), .A2(n457), .ZN(n409) );
  OR2_X1 U458 ( .A1(n670), .A2(G902), .ZN(n421) );
  XNOR2_X1 U459 ( .A(n545), .B(n447), .ZN(n678) );
  XNOR2_X1 U460 ( .A(n449), .B(n448), .ZN(n447) );
  XNOR2_X1 U461 ( .A(n531), .B(n473), .ZN(n448) );
  XNOR2_X1 U462 ( .A(n534), .B(n537), .ZN(n449) );
  NOR2_X1 U463 ( .A1(n398), .A2(n668), .ZN(n393) );
  NAND2_X1 U464 ( .A1(n401), .A2(G472), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n431), .B(n372), .ZN(n703) );
  XNOR2_X1 U466 ( .A(n682), .B(n553), .ZN(n431) );
  XNOR2_X1 U467 ( .A(G119), .B(G110), .ZN(n549) );
  INV_X1 U468 ( .A(G217), .ZN(n400) );
  XOR2_X1 U469 ( .A(KEYINPUT9), .B(G122), .Z(n521) );
  INV_X1 U470 ( .A(n659), .ZN(n596) );
  NOR2_X1 U471 ( .A1(n644), .A2(n374), .ZN(n645) );
  XNOR2_X1 U472 ( .A(G131), .B(KEYINPUT4), .ZN(n529) );
  AND2_X1 U473 ( .A1(n590), .A2(n453), .ZN(n452) );
  INV_X1 U474 ( .A(KEYINPUT45), .ZN(n453) );
  XNOR2_X1 U475 ( .A(n515), .B(n514), .ZN(n416) );
  INV_X1 U476 ( .A(KEYINPUT8), .ZN(n514) );
  XOR2_X1 U477 ( .A(G137), .B(G140), .Z(n552) );
  XOR2_X1 U478 ( .A(G107), .B(G104), .Z(n475) );
  NAND2_X1 U479 ( .A1(G234), .A2(G237), .ZN(n491) );
  NAND2_X1 U480 ( .A1(n749), .A2(n748), .ZN(n752) );
  NOR2_X1 U481 ( .A1(n760), .A2(n614), .ZN(n615) );
  BUF_X1 U482 ( .A(n569), .Z(n760) );
  XNOR2_X1 U483 ( .A(G116), .B(G101), .ZN(n535) );
  XOR2_X1 U484 ( .A(G137), .B(KEYINPUT95), .Z(n536) );
  XNOR2_X1 U485 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n532) );
  XOR2_X1 U486 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n533) );
  INV_X1 U487 ( .A(G953), .ZN(n692) );
  XNOR2_X1 U488 ( .A(n551), .B(n434), .ZN(n682) );
  INV_X1 U489 ( .A(n552), .ZN(n434) );
  XNOR2_X1 U490 ( .A(G128), .B(KEYINPUT91), .ZN(n470) );
  XNOR2_X1 U491 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n472) );
  XOR2_X1 U492 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n516) );
  XNOR2_X1 U493 ( .A(n512), .B(n511), .ZN(n670) );
  NAND2_X1 U494 ( .A1(n459), .A2(n445), .ZN(n444) );
  NAND2_X1 U495 ( .A1(n635), .A2(n461), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n387), .B(KEYINPUT41), .ZN(n777) );
  NOR2_X1 U497 ( .A1(n752), .A2(n751), .ZN(n387) );
  XOR2_X1 U498 ( .A(n500), .B(KEYINPUT0), .Z(n474) );
  BUF_X1 U499 ( .A(n764), .Z(n430) );
  NAND2_X1 U500 ( .A1(n401), .A2(G475), .ZN(n399) );
  NAND2_X1 U501 ( .A1(n401), .A2(n383), .ZN(n397) );
  NOR2_X1 U502 ( .A1(n468), .A2(n797), .ZN(n467) );
  NOR2_X1 U503 ( .A1(n796), .A2(G210), .ZN(n468) );
  NOR2_X1 U504 ( .A1(n745), .A2(n744), .ZN(n787) );
  NOR2_X1 U505 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U506 ( .A(n463), .B(n462), .ZN(n799) );
  XNOR2_X1 U507 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n462) );
  NOR2_X1 U508 ( .A1(n630), .A2(n777), .ZN(n463) );
  INV_X1 U509 ( .A(KEYINPUT40), .ZN(n464) );
  OR2_X1 U510 ( .A1(n627), .A2(n626), .ZN(n728) );
  NOR2_X1 U511 ( .A1(n629), .A2(n630), .ZN(n729) );
  XNOR2_X1 U512 ( .A(n393), .B(n384), .ZN(n679) );
  NOR2_X1 U513 ( .A1(n400), .A2(n744), .ZN(n395) );
  XNOR2_X1 U514 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U515 ( .A(n714), .B(n713), .ZN(n715) );
  AND2_X1 U516 ( .A1(n401), .A2(G469), .ZN(n369) );
  AND2_X1 U517 ( .A1(n401), .A2(G478), .ZN(n370) );
  NAND2_X1 U518 ( .A1(n488), .A2(G210), .ZN(n371) );
  XOR2_X1 U519 ( .A(n550), .B(n549), .Z(n372) );
  AND2_X1 U520 ( .A1(n435), .A2(n641), .ZN(n373) );
  OR2_X1 U521 ( .A1(n736), .A2(n643), .ZN(n374) );
  XOR2_X1 U522 ( .A(n513), .B(G475), .Z(n375) );
  NOR2_X1 U523 ( .A1(n563), .A2(n430), .ZN(n377) );
  AND2_X1 U524 ( .A1(n657), .A2(KEYINPUT48), .ZN(n378) );
  AND2_X1 U525 ( .A1(n371), .A2(n596), .ZN(n379) );
  INV_X1 U526 ( .A(n571), .ZN(n585) );
  AND2_X1 U527 ( .A1(n440), .A2(n362), .ZN(n380) );
  OR2_X1 U528 ( .A1(n371), .A2(n596), .ZN(n381) );
  INV_X1 U529 ( .A(KEYINPUT85), .ZN(n438) );
  XOR2_X1 U530 ( .A(KEYINPUT70), .B(KEYINPUT22), .Z(n382) );
  AND2_X1 U531 ( .A1(n796), .A2(G210), .ZN(n383) );
  XOR2_X1 U532 ( .A(n678), .B(KEYINPUT62), .Z(n384) );
  AND2_X1 U533 ( .A1(n577), .A2(KEYINPUT45), .ZN(n385) );
  OR2_X1 U534 ( .A1(n668), .A2(n397), .ZN(n469) );
  INV_X1 U535 ( .A(KEYINPUT44), .ZN(n455) );
  XNOR2_X2 U536 ( .A(n386), .B(n432), .ZN(n740) );
  NAND2_X1 U537 ( .A1(n386), .A2(KEYINPUT2), .ZN(n665) );
  NAND2_X2 U538 ( .A1(n414), .A2(n412), .ZN(n386) );
  NAND2_X1 U539 ( .A1(n388), .A2(n440), .ZN(n624) );
  INV_X1 U540 ( .A(n362), .ZN(n389) );
  NAND2_X1 U541 ( .A1(n396), .A2(n401), .ZN(n390) );
  NAND2_X1 U542 ( .A1(n396), .A2(n370), .ZN(n710) );
  NAND2_X1 U543 ( .A1(n396), .A2(n369), .ZN(n716) );
  NOR2_X2 U544 ( .A1(G953), .A2(n789), .ZN(n790) );
  NAND2_X1 U545 ( .A1(n391), .A2(n731), .ZN(n648) );
  XNOR2_X1 U546 ( .A(n636), .B(KEYINPUT104), .ZN(n391) );
  NAND2_X1 U547 ( .A1(n555), .A2(n554), .ZN(n392) );
  XNOR2_X1 U548 ( .A(n472), .B(KEYINPUT90), .ZN(n471) );
  INV_X1 U549 ( .A(n413), .ZN(n415) );
  NAND2_X1 U550 ( .A1(n646), .A2(n645), .ZN(n413) );
  NAND2_X2 U551 ( .A1(n444), .A2(n429), .ZN(n759) );
  NOR2_X2 U552 ( .A1(n759), .A2(n572), .ZN(n456) );
  NAND2_X1 U553 ( .A1(n407), .A2(n385), .ZN(n404) );
  XNOR2_X2 U554 ( .A(n501), .B(n474), .ZN(n571) );
  NAND2_X1 U555 ( .A1(n380), .A2(n424), .ZN(n425) );
  INV_X2 U556 ( .A(n668), .ZN(n396) );
  NAND2_X1 U557 ( .A1(n396), .A2(n395), .ZN(n704) );
  NAND2_X1 U558 ( .A1(n406), .A2(KEYINPUT45), .ZN(n405) );
  NAND2_X1 U559 ( .A1(n595), .A2(n590), .ZN(n406) );
  NAND2_X1 U560 ( .A1(n409), .A2(n408), .ZN(n411) );
  NAND2_X1 U561 ( .A1(n456), .A2(n571), .ZN(n408) );
  NAND2_X1 U562 ( .A1(n415), .A2(n378), .ZN(n414) );
  NAND2_X1 U563 ( .A1(n416), .A2(G217), .ZN(n519) );
  NAND2_X1 U564 ( .A1(n416), .A2(G221), .ZN(n553) );
  NAND2_X1 U565 ( .A1(n418), .A2(n632), .ZN(n417) );
  XNOR2_X1 U566 ( .A(n419), .B(KEYINPUT75), .ZN(n418) );
  NAND2_X1 U567 ( .A1(n628), .A2(n728), .ZN(n419) );
  XNOR2_X2 U568 ( .A(n420), .B(KEYINPUT99), .ZN(n733) );
  XNOR2_X2 U569 ( .A(n421), .B(n375), .ZN(n582) );
  INV_X1 U570 ( .A(n708), .ZN(n423) );
  NAND2_X1 U571 ( .A1(n440), .A2(n439), .ZN(n428) );
  AND2_X1 U572 ( .A1(n439), .A2(n438), .ZN(n424) );
  NAND2_X1 U573 ( .A1(n428), .A2(KEYINPUT85), .ZN(n427) );
  AND2_X2 U574 ( .A1(n427), .A2(n376), .ZN(n426) );
  AND2_X2 U575 ( .A1(n446), .A2(n460), .ZN(n429) );
  XNOR2_X1 U576 ( .A(n471), .B(n470), .ZN(n550) );
  NAND2_X1 U577 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U578 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X2 U579 ( .A(n683), .B(G146), .ZN(n545) );
  NOR2_X2 U580 ( .A1(G902), .A2(n712), .ZN(n548) );
  INV_X1 U581 ( .A(n734), .ZN(n437) );
  NAND2_X1 U582 ( .A1(n442), .A2(KEYINPUT66), .ZN(n594) );
  NAND2_X1 U583 ( .A1(n443), .A2(n455), .ZN(n442) );
  XNOR2_X1 U584 ( .A(n591), .B(KEYINPUT68), .ZN(n443) );
  AND2_X1 U585 ( .A1(n657), .A2(n647), .ZN(n450) );
  XNOR2_X2 U586 ( .A(n451), .B(n382), .ZN(n539) );
  XNOR2_X2 U587 ( .A(n565), .B(n564), .ZN(n676) );
  XNOR2_X2 U588 ( .A(G143), .B(G128), .ZN(n520) );
  NAND2_X1 U589 ( .A1(n585), .A2(n572), .ZN(n458) );
  NAND2_X1 U590 ( .A1(n759), .A2(n572), .ZN(n457) );
  NAND2_X1 U591 ( .A1(n586), .A2(n461), .ZN(n460) );
  INV_X1 U592 ( .A(KEYINPUT33), .ZN(n461) );
  NAND2_X1 U593 ( .A1(n655), .A2(n633), .ZN(n465) );
  XNOR2_X1 U594 ( .A(n611), .B(n610), .ZN(n655) );
  NAND2_X1 U595 ( .A1(n469), .A2(n467), .ZN(n466) );
  AND2_X1 U596 ( .A1(n530), .A2(G210), .ZN(n473) );
  XNOR2_X1 U597 ( .A(n552), .B(n475), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n677), .A2(n656), .ZN(n657) );
  XNOR2_X1 U599 ( .A(n551), .B(n507), .ZN(n512) );
  XNOR2_X2 U600 ( .A(G110), .B(G101), .ZN(n540) );
  XNOR2_X2 U601 ( .A(G116), .B(G107), .ZN(n517) );
  XNOR2_X1 U602 ( .A(n540), .B(n517), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n503), .B(KEYINPUT16), .ZN(n476) );
  XNOR2_X1 U604 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U605 ( .A(KEYINPUT3), .B(G119), .ZN(n478) );
  XNOR2_X1 U606 ( .A(n478), .B(G113), .ZN(n531) );
  XNOR2_X2 U607 ( .A(n480), .B(G953), .ZN(n684) );
  NAND2_X1 U608 ( .A1(n684), .A2(G224), .ZN(n483) );
  XNOR2_X1 U609 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n481) );
  XNOR2_X1 U610 ( .A(n481), .B(KEYINPUT4), .ZN(n482) );
  XNOR2_X1 U611 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X2 U612 ( .A(G125), .B(G146), .ZN(n506) );
  XNOR2_X1 U613 ( .A(n520), .B(n506), .ZN(n484) );
  XNOR2_X1 U614 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U615 ( .A(KEYINPUT15), .B(G902), .ZN(n659) );
  XNOR2_X1 U616 ( .A(KEYINPUT71), .B(n487), .ZN(n488) );
  NAND2_X1 U617 ( .A1(n488), .A2(G214), .ZN(n490) );
  INV_X1 U618 ( .A(KEYINPUT87), .ZN(n489) );
  XNOR2_X1 U619 ( .A(n490), .B(n489), .ZN(n748) );
  INV_X1 U620 ( .A(n748), .ZN(n651) );
  XNOR2_X1 U621 ( .A(n491), .B(KEYINPUT14), .ZN(n747) );
  AND2_X1 U622 ( .A1(n692), .A2(G952), .ZN(n492) );
  AND2_X1 U623 ( .A1(n747), .A2(n492), .ZN(n601) );
  INV_X1 U624 ( .A(n601), .ZN(n498) );
  INV_X1 U625 ( .A(G898), .ZN(n493) );
  NAND2_X1 U626 ( .A1(n493), .A2(G953), .ZN(n495) );
  INV_X1 U627 ( .A(KEYINPUT88), .ZN(n494) );
  XNOR2_X1 U628 ( .A(n495), .B(n494), .ZN(n699) );
  AND2_X1 U629 ( .A1(n699), .A2(G902), .ZN(n496) );
  NAND2_X1 U630 ( .A1(n496), .A2(n747), .ZN(n497) );
  AND2_X1 U631 ( .A1(n498), .A2(n497), .ZN(n499) );
  INV_X1 U632 ( .A(KEYINPUT86), .ZN(n500) );
  XNOR2_X1 U633 ( .A(n363), .B(n502), .ZN(n505) );
  XNOR2_X1 U634 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U635 ( .A(n506), .B(KEYINPUT10), .ZN(n551) );
  NAND2_X1 U636 ( .A1(G214), .A2(n530), .ZN(n509) );
  XNOR2_X1 U637 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U638 ( .A(n510), .B(KEYINPUT96), .Z(n511) );
  XNOR2_X1 U639 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n513) );
  NAND2_X1 U640 ( .A1(n684), .A2(G234), .ZN(n515) );
  XNOR2_X1 U641 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U642 ( .A(n519), .B(n518), .ZN(n523) );
  XNOR2_X1 U643 ( .A(n528), .B(n521), .ZN(n522) );
  XNOR2_X1 U644 ( .A(n523), .B(n522), .ZN(n708) );
  INV_X1 U645 ( .A(n583), .ZN(n573) );
  AND2_X1 U646 ( .A1(n582), .A2(n573), .ZN(n613) );
  NAND2_X1 U647 ( .A1(G234), .A2(n659), .ZN(n524) );
  XNOR2_X1 U648 ( .A(KEYINPUT20), .B(n524), .ZN(n556) );
  NAND2_X1 U649 ( .A1(n556), .A2(G221), .ZN(n526) );
  INV_X1 U650 ( .A(KEYINPUT21), .ZN(n525) );
  XNOR2_X1 U651 ( .A(n526), .B(n525), .ZN(n761) );
  AND2_X1 U652 ( .A1(n613), .A2(n761), .ZN(n527) );
  XNOR2_X1 U653 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U654 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U655 ( .A1(n678), .A2(n554), .ZN(n538) );
  XNOR2_X1 U656 ( .A(n540), .B(KEYINPUT89), .ZN(n542) );
  NAND2_X1 U657 ( .A1(n684), .A2(G227), .ZN(n541) );
  XNOR2_X1 U658 ( .A(n542), .B(n541), .ZN(n544) );
  INV_X1 U659 ( .A(G469), .ZN(n547) );
  XNOR2_X2 U660 ( .A(n548), .B(n547), .ZN(n620) );
  XNOR2_X2 U661 ( .A(n620), .B(KEYINPUT1), .ZN(n649) );
  INV_X1 U662 ( .A(n703), .ZN(n555) );
  INV_X1 U663 ( .A(G902), .ZN(n554) );
  NAND2_X1 U664 ( .A1(n556), .A2(G217), .ZN(n558) );
  XNOR2_X1 U665 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n557) );
  INV_X1 U666 ( .A(n760), .ZN(n579) );
  AND2_X1 U667 ( .A1(n649), .A2(n579), .ZN(n560) );
  INV_X1 U668 ( .A(KEYINPUT32), .ZN(n561) );
  OR2_X1 U669 ( .A1(n649), .A2(n760), .ZN(n563) );
  INV_X1 U670 ( .A(KEYINPUT101), .ZN(n564) );
  NAND2_X1 U671 ( .A1(n676), .A2(KEYINPUT68), .ZN(n566) );
  NOR2_X1 U672 ( .A1(n681), .A2(n566), .ZN(n567) );
  INV_X1 U673 ( .A(n567), .ZN(n568) );
  NAND2_X1 U674 ( .A1(n568), .A2(KEYINPUT66), .ZN(n576) );
  INV_X1 U675 ( .A(n766), .ZN(n570) );
  INV_X1 U676 ( .A(KEYINPUT34), .ZN(n572) );
  AND2_X1 U677 ( .A1(n365), .A2(KEYINPUT44), .ZN(n575) );
  NAND2_X1 U678 ( .A1(n455), .A2(KEYINPUT66), .ZN(n577) );
  INV_X1 U679 ( .A(KEYINPUT84), .ZN(n578) );
  XNOR2_X1 U680 ( .A(n366), .B(n578), .ZN(n581) );
  NOR2_X1 U681 ( .A1(n649), .A2(n579), .ZN(n580) );
  AND2_X1 U682 ( .A1(n581), .A2(n580), .ZN(n718) );
  NOR2_X1 U683 ( .A1(n583), .A2(n582), .ZN(n633) );
  NOR2_X1 U684 ( .A1(n733), .A2(n633), .ZN(n584) );
  XNOR2_X1 U685 ( .A(n584), .B(KEYINPUT100), .ZN(n753) );
  INV_X1 U686 ( .A(n753), .ZN(n641) );
  INV_X1 U687 ( .A(n430), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n586), .A2(n616), .ZN(n773) );
  NAND2_X1 U689 ( .A1(n571), .A2(n773), .ZN(n587) );
  XNOR2_X1 U690 ( .A(n587), .B(KEYINPUT31), .ZN(n734) );
  INV_X1 U691 ( .A(n766), .ZN(n588) );
  NAND2_X1 U692 ( .A1(n588), .A2(n620), .ZN(n604) );
  NOR2_X1 U693 ( .A1(n430), .A2(n604), .ZN(n589) );
  AND2_X1 U694 ( .A1(n571), .A2(n589), .ZN(n721) );
  INV_X1 U695 ( .A(n681), .ZN(n592) );
  AND2_X1 U696 ( .A1(n592), .A2(n676), .ZN(n593) );
  NAND2_X1 U697 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U698 ( .A1(n666), .A2(n596), .ZN(n597) );
  XNOR2_X1 U699 ( .A(n597), .B(KEYINPUT79), .ZN(n658) );
  NAND2_X1 U700 ( .A1(G902), .A2(n747), .ZN(n598) );
  NOR2_X1 U701 ( .A1(G900), .A2(n598), .ZN(n599) );
  INV_X1 U702 ( .A(n684), .ZN(n672) );
  NAND2_X1 U703 ( .A1(n599), .A2(n672), .ZN(n600) );
  XNOR2_X1 U704 ( .A(n600), .B(KEYINPUT103), .ZN(n602) );
  NOR2_X1 U705 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U706 ( .A(KEYINPUT74), .B(n603), .ZN(n614) );
  XNOR2_X1 U707 ( .A(n605), .B(KEYINPUT72), .ZN(n609) );
  NAND2_X1 U708 ( .A1(n748), .A2(n764), .ZN(n606) );
  XNOR2_X1 U709 ( .A(n606), .B(KEYINPUT30), .ZN(n607) );
  XNOR2_X1 U710 ( .A(KEYINPUT105), .B(n607), .ZN(n608) );
  NAND2_X1 U711 ( .A1(n609), .A2(n608), .ZN(n627) );
  XNOR2_X1 U712 ( .A(KEYINPUT69), .B(KEYINPUT39), .ZN(n610) );
  INV_X1 U713 ( .A(n613), .ZN(n751) );
  NAND2_X1 U714 ( .A1(n615), .A2(n761), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n617) );
  XNOR2_X1 U716 ( .A(KEYINPUT28), .B(n617), .ZN(n618) );
  XNOR2_X1 U717 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U718 ( .A1(n621), .A2(n620), .ZN(n630) );
  XNOR2_X1 U719 ( .A(n622), .B(KEYINPUT46), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n753), .A2(KEYINPUT47), .ZN(n623) );
  XNOR2_X1 U721 ( .A(n623), .B(KEYINPUT78), .ZN(n628) );
  INV_X1 U722 ( .A(n624), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n625), .A2(n653), .ZN(n626) );
  INV_X1 U724 ( .A(n729), .ZN(n631) );
  NAND2_X1 U725 ( .A1(n631), .A2(KEYINPUT47), .ZN(n632) );
  INV_X1 U726 ( .A(n649), .ZN(n767) );
  XNOR2_X1 U727 ( .A(KEYINPUT102), .B(n633), .ZN(n731) );
  NOR2_X1 U728 ( .A1(n635), .A2(n634), .ZN(n636) );
  INV_X1 U729 ( .A(n648), .ZN(n638) );
  NAND2_X1 U730 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U731 ( .A(n639), .B(KEYINPUT36), .ZN(n640) );
  NOR2_X1 U732 ( .A1(n767), .A2(n640), .ZN(n736) );
  NAND2_X1 U733 ( .A1(n641), .A2(n729), .ZN(n642) );
  NOR2_X1 U734 ( .A1(KEYINPUT47), .A2(n642), .ZN(n643) );
  INV_X1 U735 ( .A(KEYINPUT48), .ZN(n647) );
  OR2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U737 ( .A(n652), .B(KEYINPUT43), .ZN(n654) );
  NOR2_X1 U738 ( .A1(n654), .A2(n653), .ZN(n677) );
  NAND2_X1 U739 ( .A1(n733), .A2(n655), .ZN(n739) );
  NAND2_X1 U740 ( .A1(n658), .A2(n740), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT80), .B(n659), .Z(n660) );
  NAND2_X1 U742 ( .A1(n660), .A2(KEYINPUT2), .ZN(n661) );
  XNOR2_X2 U743 ( .A(n664), .B(KEYINPUT65), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n665), .B(KEYINPUT82), .ZN(n667) );
  INV_X1 U745 ( .A(n360), .ZN(n741) );
  XOR2_X1 U746 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n669) );
  INV_X1 U747 ( .A(G952), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n705) );
  NAND2_X1 U749 ( .A1(n673), .A2(n705), .ZN(n675) );
  INV_X1 U750 ( .A(KEYINPUT60), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n675), .B(n674), .ZN(G60) );
  XNOR2_X1 U752 ( .A(n676), .B(G110), .ZN(G12) );
  XNOR2_X1 U753 ( .A(n365), .B(G122), .ZN(G24) );
  XOR2_X1 U754 ( .A(n677), .B(G140), .Z(G42) );
  NAND2_X1 U755 ( .A1(n679), .A2(n705), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n680), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U757 ( .A(n681), .B(G119), .Z(G21) );
  XOR2_X1 U758 ( .A(n683), .B(n682), .Z(n686) );
  XOR2_X1 U759 ( .A(n686), .B(n740), .Z(n685) );
  NAND2_X1 U760 ( .A1(n685), .A2(n684), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n686), .B(G227), .ZN(n687) );
  XNOR2_X1 U762 ( .A(n687), .B(KEYINPUT126), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n688), .A2(G900), .ZN(n689) );
  NAND2_X1 U764 ( .A1(G953), .A2(n689), .ZN(n690) );
  NAND2_X1 U765 ( .A1(n691), .A2(n690), .ZN(G72) );
  NAND2_X1 U766 ( .A1(n360), .A2(n692), .ZN(n697) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n693) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n693), .ZN(n694) );
  NAND2_X1 U769 ( .A1(n694), .A2(G898), .ZN(n695) );
  XNOR2_X1 U770 ( .A(n695), .B(KEYINPUT124), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n697), .A2(n696), .ZN(n702) );
  NOR2_X1 U772 ( .A1(n698), .A2(n699), .ZN(n700) );
  XOR2_X1 U773 ( .A(KEYINPUT125), .B(n700), .Z(n701) );
  XNOR2_X1 U774 ( .A(n702), .B(n701), .ZN(G69) );
  XNOR2_X1 U775 ( .A(n703), .B(n704), .ZN(n706) );
  INV_X1 U776 ( .A(n705), .ZN(n797) );
  NOR2_X1 U777 ( .A1(n706), .A2(n797), .ZN(G66) );
  XOR2_X1 U778 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n707) );
  XNOR2_X1 U779 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n711), .A2(n797), .ZN(G63) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n714) );
  XNOR2_X1 U782 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  XNOR2_X1 U783 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n717), .A2(n797), .ZN(G54) );
  XNOR2_X1 U785 ( .A(G101), .B(n718), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U787 ( .A1(n731), .A2(n721), .ZN(n720) );
  XNOR2_X1 U788 ( .A(n720), .B(G104), .ZN(G6) );
  XNOR2_X1 U789 ( .A(G107), .B(KEYINPUT27), .ZN(n725) );
  XOR2_X1 U790 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n723) );
  NAND2_X1 U791 ( .A1(n721), .A2(n733), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U793 ( .A(n725), .B(n724), .ZN(G9) );
  XOR2_X1 U794 ( .A(G128), .B(KEYINPUT29), .Z(n727) );
  NAND2_X1 U795 ( .A1(n729), .A2(n733), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n727), .B(n726), .ZN(G30) );
  XNOR2_X1 U797 ( .A(G143), .B(n728), .ZN(G45) );
  NAND2_X1 U798 ( .A1(n729), .A2(n731), .ZN(n730) );
  XNOR2_X1 U799 ( .A(n730), .B(G146), .ZN(G48) );
  NAND2_X1 U800 ( .A1(n731), .A2(n734), .ZN(n732) );
  XNOR2_X1 U801 ( .A(n732), .B(G113), .ZN(G15) );
  NAND2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U803 ( .A(n735), .B(G116), .ZN(G18) );
  XNOR2_X1 U804 ( .A(G125), .B(n736), .ZN(n737) );
  XNOR2_X1 U805 ( .A(n737), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U806 ( .A(G134), .B(KEYINPUT111), .Z(n738) );
  XNOR2_X1 U807 ( .A(n739), .B(n738), .ZN(G36) );
  INV_X1 U808 ( .A(n740), .ZN(n742) );
  NOR2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U810 ( .A1(n743), .A2(KEYINPUT2), .ZN(n745) );
  NOR2_X1 U811 ( .A1(n759), .A2(n777), .ZN(n746) );
  XNOR2_X1 U812 ( .A(n746), .B(KEYINPUT117), .ZN(n785) );
  INV_X1 U813 ( .A(n747), .ZN(n782) );
  NOR2_X1 U814 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U815 ( .A1(n751), .A2(n750), .ZN(n756) );
  NOR2_X1 U816 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U817 ( .A(KEYINPUT115), .B(n754), .Z(n755) );
  NOR2_X1 U818 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U819 ( .A(n757), .B(KEYINPUT116), .ZN(n758) );
  NOR2_X1 U820 ( .A1(n759), .A2(n758), .ZN(n779) );
  NOR2_X1 U821 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U822 ( .A(KEYINPUT49), .B(n762), .Z(n763) );
  NOR2_X1 U823 ( .A1(n430), .A2(n763), .ZN(n765) );
  XOR2_X1 U824 ( .A(KEYINPUT112), .B(n765), .Z(n771) );
  NAND2_X1 U825 ( .A1(n766), .A2(n767), .ZN(n768) );
  XNOR2_X1 U826 ( .A(n768), .B(KEYINPUT113), .ZN(n769) );
  XNOR2_X1 U827 ( .A(KEYINPUT50), .B(n769), .ZN(n770) );
  NOR2_X1 U828 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U829 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U830 ( .A(KEYINPUT51), .B(n774), .Z(n775) );
  XNOR2_X1 U831 ( .A(n775), .B(KEYINPUT114), .ZN(n776) );
  NOR2_X1 U832 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U833 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U834 ( .A(n780), .B(KEYINPUT52), .ZN(n781) );
  NOR2_X1 U835 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U836 ( .A1(n783), .A2(G952), .ZN(n784) );
  NAND2_X1 U837 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U838 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U839 ( .A(KEYINPUT118), .B(n788), .Z(n789) );
  XNOR2_X1 U840 ( .A(KEYINPUT53), .B(n790), .ZN(G75) );
  XOR2_X1 U841 ( .A(KEYINPUT55), .B(KEYINPUT76), .Z(n792) );
  XNOR2_X1 U842 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n791) );
  XNOR2_X1 U843 ( .A(n792), .B(n791), .ZN(n794) );
  XOR2_X1 U844 ( .A(n794), .B(n793), .Z(n795) );
  INV_X1 U845 ( .A(n795), .ZN(n796) );
  XNOR2_X1 U846 ( .A(n798), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U847 ( .A(G137), .B(n799), .ZN(n800) );
  XNOR2_X1 U848 ( .A(n800), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U849 ( .A(n801), .B(G131), .Z(G33) );
endmodule

