//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT66), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n207), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n228), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n216), .A2(new_n217), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n220), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n256), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n219), .A2(new_n256), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n267), .B2(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G159), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n255), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT81), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n229), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n259), .A2(new_n265), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n271), .B1(new_n278), .B2(G68), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n279), .B2(KEYINPUT16), .ZN(new_n280));
  OAI211_X1 g0080(.A(KEYINPUT81), .B(new_n255), .C1(new_n266), .C2(new_n271), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n229), .A3(new_n275), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n219), .A2(KEYINPUT8), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n285), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n261), .A2(new_n263), .A3(G223), .A4(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(G33), .A2(G41), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n229), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  INV_X1    g0110(.A(G45), .ZN(new_n311));
  AOI21_X1  g0111(.A(G1), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G274), .ZN(new_n314));
  AND2_X1   g0114(.A1(G1), .A2(G13), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n313), .A2(G232), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n309), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n309), .A2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(G200), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n282), .A2(new_n301), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT17), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n282), .A2(KEYINPUT17), .A3(new_n301), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n261), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(new_n302), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n308), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n313), .A2(G238), .B1(new_n312), .B2(new_n317), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n332), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g0136(.A(G200), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n333), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(G190), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n269), .A2(G50), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n230), .A2(G33), .A3(G77), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n256), .A2(G20), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT11), .B1(new_n345), .B2(new_n276), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT76), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n276), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT11), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT76), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n346), .ZN(new_n354));
  INV_X1    g0154(.A(new_n286), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n284), .A2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT77), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n286), .B2(new_n356), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n358), .A2(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n349), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n337), .A2(new_n341), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT78), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n337), .A2(new_n341), .A3(new_n364), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n349), .A2(new_n354), .A3(new_n363), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n335), .A2(new_n336), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n373));
  OAI211_X1 g0173(.A(G169), .B(new_n373), .C1(new_n335), .C2(new_n336), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n339), .A2(new_n340), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(G169), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n282), .A2(new_n301), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n309), .A2(new_n318), .A3(G179), .ZN(new_n381));
  INV_X1    g0181(.A(G169), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n309), .B2(new_n318), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT82), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n282), .B2(new_n301), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n380), .B2(new_n385), .ZN(new_n393));
  AOI211_X1 g0193(.A(KEYINPUT18), .B(new_n384), .C1(new_n282), .C2(new_n301), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT82), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI211_X1 g0195(.A(new_n327), .B(new_n379), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n230), .A2(G33), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n294), .A2(new_n297), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n203), .A2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n203), .A2(KEYINPUT71), .A3(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n269), .A2(G150), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n276), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(G50), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n300), .A2(new_n202), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n317), .A2(new_n312), .ZN(new_n410));
  INV_X1    g0210(.A(G226), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n316), .A2(G1), .A3(G13), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n410), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n258), .A2(G222), .A3(new_n302), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n264), .A2(G77), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n419), .B2(new_n308), .ZN(new_n420));
  INV_X1    g0220(.A(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n409), .B(new_n422), .C1(G169), .C2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n300), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n284), .A2(G77), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n286), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n293), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n397), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n430), .B2(new_n276), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n258), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n264), .A2(new_n220), .A3(G1698), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n308), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G244), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n410), .B1(new_n437), .B2(new_n414), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT73), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n410), .B(KEYINPUT73), .C1(new_n437), .C2(new_n414), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n431), .B1(new_n442), .B2(new_n382), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n436), .A2(new_n421), .A3(new_n440), .A4(new_n441), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(G200), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n436), .A2(G190), .A3(new_n440), .A4(new_n441), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n431), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n420), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n419), .A2(new_n308), .ZN(new_n453));
  INV_X1    g0253(.A(new_n415), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT74), .A3(G200), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT9), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n409), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT9), .A4(new_n408), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n420), .A2(G190), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n460), .A2(KEYINPUT10), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT10), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n452), .A2(new_n456), .B1(new_n409), .B2(new_n458), .ZN(new_n466));
  INV_X1    g0266(.A(new_n463), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n423), .B(new_n449), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT75), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT10), .B1(new_n460), .B2(new_n463), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n467), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT75), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n423), .A4(new_n449), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n396), .A2(new_n476), .A3(KEYINPUT83), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT83), .B1(new_n396), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n261), .A2(new_n263), .A3(new_n230), .A4(G87), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n258), .A2(new_n230), .A3(G87), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n230), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n433), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n482), .A2(new_n485), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n277), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n285), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n283), .A2(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n285), .A2(new_n499), .A3(new_n229), .A4(new_n275), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n433), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n261), .A2(new_n263), .A3(G257), .A4(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(new_n302), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n308), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n311), .A2(G1), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT5), .B(G41), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n317), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n508), .B1(new_n315), .B2(new_n316), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G264), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n506), .A2(new_n308), .B1(new_n511), .B2(G264), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT90), .A3(new_n510), .ZN(new_n517));
  AOI21_X1  g0317(.A(G190), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n513), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G200), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n502), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n510), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(G257), .B2(new_n511), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(new_n302), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(KEYINPUT85), .A3(new_n527), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n523), .B1(new_n533), .B2(new_n412), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(KEYINPUT6), .B2(new_n221), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(G20), .C1(new_n536), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n269), .A2(G77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n433), .B1(new_n259), .B2(new_n265), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n276), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n300), .A2(new_n221), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n500), .B2(new_n221), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G190), .B(new_n523), .C1(new_n533), .C2(new_n412), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n535), .A2(new_n545), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n355), .A2(new_n551), .A3(G87), .A4(new_n499), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT87), .B1(new_n500), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n221), .A3(new_n433), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(new_n221), .A3(new_n433), .A4(KEYINPUT86), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(new_n559), .B1(new_n230), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n261), .A2(new_n263), .A3(new_n230), .A4(G68), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n397), .A2(new_n221), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(KEYINPUT19), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n276), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n429), .A2(new_n300), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n412), .A2(G274), .A3(new_n508), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n283), .A2(G45), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(G250), .C1(new_n307), .C2(new_n229), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n261), .A2(new_n263), .A3(G238), .A4(new_n302), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(new_n486), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n319), .B(new_n571), .C1(new_n308), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n574), .B2(new_n308), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  AOI211_X1 g0379(.A(G179), .B(new_n571), .C1(new_n308), .C2(new_n574), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n308), .ZN(new_n581));
  INV_X1    g0381(.A(new_n571), .ZN(new_n582));
  AOI21_X1  g0382(.A(G169), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n565), .B(new_n566), .C1(new_n429), .C2(new_n500), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n576), .A2(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n545), .A2(new_n548), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n421), .B(new_n523), .C1(new_n533), .C2(new_n412), .ZN(new_n588));
  INV_X1    g0388(.A(new_n511), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n510), .B1(new_n589), .B2(new_n222), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n526), .A2(new_n527), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n525), .A2(new_n524), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n526), .A2(KEYINPUT85), .A3(new_n527), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT85), .B1(new_n526), .B2(new_n527), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n590), .B1(new_n595), .B2(new_n308), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n587), .B(new_n588), .C1(G169), .C2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n521), .A2(new_n550), .A3(new_n586), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n515), .A2(G169), .A3(new_n517), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n519), .A2(G179), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT91), .ZN(new_n602));
  INV_X1    g0402(.A(new_n502), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n264), .A2(G303), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n261), .A2(new_n263), .A3(G264), .A4(G1698), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n261), .A2(new_n263), .A3(G257), .A4(new_n302), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(KEYINPUT88), .A3(new_n609), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n308), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n524), .B(new_n230), .C1(G33), .C2(new_n221), .ZN(new_n617));
  INV_X1    g0417(.A(G116), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G20), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n276), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n620), .B(new_n621), .ZN(new_n622));
  MUX2_X1   g0422(.A(new_n285), .B(new_n500), .S(G116), .Z(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(KEYINPUT5), .A2(G41), .ZN(new_n625));
  NOR2_X1   g0425(.A1(KEYINPUT5), .A2(G41), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n508), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(G270), .A3(new_n412), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n628), .A2(G179), .A3(new_n510), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n616), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n412), .B1(new_n613), .B2(new_n614), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n510), .ZN(new_n633));
  OAI211_X1 g0433(.A(G169), .B(new_n624), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT21), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n382), .B1(new_n622), .B2(new_n623), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n633), .C2(new_n632), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n631), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n624), .ZN(new_n640));
  OAI21_X1  g0440(.A(G200), .B1(new_n632), .B2(new_n633), .ZN(new_n641));
  INV_X1    g0441(.A(new_n633), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n616), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n641), .C1(new_n643), .C2(new_n319), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n479), .A2(new_n598), .A3(new_n607), .A4(new_n645), .ZN(G372));
  AND3_X1   g0446(.A1(new_n443), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT92), .B1(new_n443), .B2(new_n444), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n365), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n327), .B1(new_n650), .B2(new_n378), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n393), .A2(new_n394), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n473), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n423), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n597), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n586), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n584), .A2(new_n585), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n565), .A2(new_n566), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n577), .A2(G190), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n579), .A2(new_n661), .A3(new_n555), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n659), .B1(new_n664), .B2(new_n597), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n601), .A2(new_n603), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n598), .B1(new_n668), .B2(new_n639), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n656), .B1(new_n479), .B2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n635), .A2(new_n638), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n630), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n283), .A2(new_n230), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT93), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n601), .A2(new_n603), .A3(new_n679), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n521), .B1(new_n502), .B2(new_n680), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n607), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n502), .B1(new_n599), .B2(new_n600), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n682), .A2(new_n685), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n640), .A2(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n645), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n212), .A2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n233), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n558), .A2(new_n618), .A3(new_n559), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G1), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n597), .A2(new_n521), .A3(new_n550), .A4(new_n586), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n686), .B2(new_n673), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n658), .A2(new_n665), .B1(new_n585), .B2(new_n584), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n679), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n668), .A2(KEYINPUT91), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n686), .A2(new_n602), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n639), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n700), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n679), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n705), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n516), .A2(new_n629), .A3(new_n577), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n596), .A2(new_n712), .A3(new_n616), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n596), .A2(new_n712), .A3(KEYINPUT30), .A4(new_n616), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n578), .A2(new_n513), .A3(new_n421), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n643), .A2(new_n717), .A3(new_n534), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n719), .B2(new_n679), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n672), .A2(new_n630), .A3(new_n644), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n606), .A2(new_n700), .A3(new_n723), .A4(new_n680), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n711), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n699), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(G13), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n283), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n694), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n691), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G330), .B2(new_n690), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n315), .B1(new_n230), .B2(G169), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n249), .A2(new_n311), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n212), .A2(new_n258), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n745), .B(new_n747), .C1(new_n311), .C2(new_n233), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n213), .A2(G355), .A3(new_n258), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G116), .B2(new_n213), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n744), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n734), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n319), .A2(G20), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT97), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n421), .A2(new_n451), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G329), .ZN(new_n762));
  NAND2_X1  g0562(.A1(G20), .A2(G179), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n451), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(new_n319), .A3(new_n451), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G326), .A2(new_n766), .B1(new_n768), .B2(G311), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(G190), .A3(new_n451), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n764), .A2(new_n319), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G322), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  OAI21_X1  g0576(.A(G20), .B1(new_n756), .B2(new_n319), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n421), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n264), .B1(new_n776), .B2(new_n778), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n755), .A2(G179), .A3(new_n451), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G283), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n762), .A2(new_n769), .A3(new_n775), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n761), .A2(G159), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n790), .A2(new_n202), .B1(new_n424), .B2(new_n767), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G68), .B2(new_n773), .ZN(new_n792));
  INV_X1    g0592(.A(new_n782), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G87), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n777), .A2(G97), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n258), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G107), .B2(new_n785), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n770), .B(KEYINPUT96), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n792), .B(new_n797), .C1(new_n219), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n787), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n752), .B1(new_n740), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n743), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n690), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n736), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n648), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n443), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n431), .A2(new_n680), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n808), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n445), .A2(new_n448), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n703), .B(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n734), .B1(new_n813), .B2(new_n726), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n726), .B2(new_n813), .ZN(new_n815));
  INV_X1    g0615(.A(new_n740), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n258), .B1(new_n778), .B2(new_n219), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G68), .B2(new_n785), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n202), .B2(new_n782), .C1(new_n760), .C2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G137), .A2(new_n766), .B1(new_n768), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  INV_X1    g0622(.A(G143), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n822), .B2(new_n772), .C1(new_n798), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT101), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n761), .A2(G311), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n785), .A2(G87), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n264), .A3(new_n795), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G107), .B2(new_n793), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G303), .A2(new_n766), .B1(new_n773), .B2(G283), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G116), .A2(new_n768), .B1(new_n771), .B2(G294), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n829), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n816), .B1(new_n836), .B2(KEYINPUT102), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT102), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n740), .A2(new_n741), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n734), .B1(G77), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  OAI211_X1 g0642(.A(new_n838), .B(new_n842), .C1(new_n742), .C2(new_n812), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n815), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  OAI21_X1  g0645(.A(new_n539), .B1(new_n536), .B2(new_n540), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT35), .ZN(new_n847));
  OAI211_X1 g0647(.A(G116), .B(new_n231), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT36), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n233), .B(G77), .C1(new_n219), .C2(new_n256), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n202), .A2(G68), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n283), .B(G13), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n677), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n380), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n386), .A2(new_n856), .A3(new_n857), .A4(new_n323), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n280), .A2(new_n272), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n301), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n385), .B2(new_n855), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n861), .A2(new_n323), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n858), .B1(new_n862), .B2(new_n857), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n327), .B1(new_n392), .B2(new_n395), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n855), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n370), .A2(new_n679), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n375), .A2(new_n377), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n369), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n365), .A2(new_n871), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT79), .B(KEYINPUT14), .C1(new_n371), .C2(new_n382), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n372), .A3(new_n374), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n876), .B2(new_n370), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n812), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n724), .B2(new_n722), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT40), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n445), .A2(new_n448), .A3(new_n810), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n649), .B2(new_n808), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n370), .B1(new_n371), .B2(G190), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n367), .B1(new_n883), .B2(new_n337), .ZN(new_n884));
  INV_X1    g0684(.A(new_n368), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n871), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n877), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n725), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n869), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n282), .A2(new_n301), .A3(new_n322), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n389), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n857), .B1(new_n896), .B2(new_n856), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n387), .A2(new_n325), .A3(new_n326), .A4(new_n391), .ZN(new_n898));
  INV_X1    g0698(.A(new_n856), .ZN(new_n899));
  AOI22_X1  g0699(.A1(KEYINPUT104), .A2(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n386), .A2(new_n856), .A3(new_n323), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n858), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n893), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT40), .B1(new_n891), .B2(new_n892), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT106), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n898), .A2(new_n899), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n867), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n912), .A2(new_n869), .B1(new_n891), .B2(new_n892), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT106), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n879), .B2(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n880), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n479), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n918), .A2(new_n919), .A3(new_n725), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n725), .ZN(new_n921));
  INV_X1    g0721(.A(G330), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT107), .Z(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n894), .B2(new_n905), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n876), .A2(new_n370), .A3(new_n680), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n888), .A2(new_n889), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n680), .B(new_n812), .C1(new_n667), .C2(new_n669), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n443), .A2(new_n444), .A3(new_n680), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT103), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n932), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n870), .A2(new_n937), .B1(new_n653), .B2(new_n677), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n711), .B1(new_n477), .B2(new_n478), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n656), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n939), .B(new_n941), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n924), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(G1), .B1(new_n730), .B2(G20), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(KEYINPUT108), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n924), .B2(new_n942), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT108), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n854), .B1(new_n946), .B2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n567), .A2(new_n679), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n586), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n660), .A2(new_n949), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n587), .A2(new_n679), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n550), .A2(new_n597), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n597), .B2(new_n680), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n682), .A2(new_n685), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n606), .A2(new_n958), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n679), .B1(new_n962), .B2(new_n597), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n956), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n954), .A2(new_n955), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n692), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n959), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n967), .B(new_n969), .Z(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n694), .B(new_n971), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n687), .A2(new_n959), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT111), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n687), .A2(new_n976), .A3(new_n959), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n687), .A2(new_n959), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(new_n968), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n691), .A2(new_n685), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n692), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n682), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n968), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n728), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n973), .B1(new_n990), .B2(new_n728), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n970), .B1(new_n991), .B2(new_n733), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n782), .A2(new_n618), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(KEYINPUT46), .B1(new_n768), .B2(G283), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n766), .B1(new_n773), .B2(G294), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n785), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n221), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n258), .B(new_n998), .C1(G107), .C2(new_n777), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(KEYINPUT46), .B2(new_n993), .C1(new_n1000), .C2(new_n760), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n798), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n996), .B(new_n1001), .C1(G303), .C2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n761), .A2(G137), .B1(G58), .B2(new_n793), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n785), .A2(G77), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n778), .A2(new_n256), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n264), .ZN(new_n1010));
  INV_X1    g0810(.A(G159), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1008), .B(new_n1010), .C1(new_n1011), .C2(new_n772), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G143), .A2(new_n766), .B1(new_n771), .B2(G150), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n202), .B2(new_n767), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1007), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1003), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n816), .B1(new_n1016), .B2(KEYINPUT47), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT47), .B2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n954), .A2(new_n743), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n734), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n746), .A2(new_n239), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n429), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n743), .B(new_n740), .C1(new_n212), .C2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n992), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT113), .ZN(G387));
  INV_X1    g0827(.A(new_n694), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n988), .B2(new_n728), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n728), .B2(new_n988), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n244), .A2(G45), .A3(new_n264), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT50), .B1(new_n295), .B2(G50), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n311), .C1(new_n256), .C2(new_n424), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n295), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n264), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n696), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n212), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n744), .B1(new_n213), .B2(new_n433), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n768), .B1(new_n773), .B2(new_n298), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n202), .B2(new_n770), .C1(new_n1011), .C2(new_n790), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n782), .A2(new_n424), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n778), .A2(new_n429), .ZN(new_n1042));
  OR4_X1    g0842(.A1(new_n264), .A2(new_n998), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G150), .C2(new_n761), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G303), .A2(new_n768), .B1(new_n773), .B2(G311), .ZN(new_n1045));
  INV_X1    g0845(.A(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n790), .C1(new_n798), .C2(new_n1000), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n793), .A2(G294), .B1(G283), .B2(new_n777), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n264), .B1(new_n997), .B2(new_n618), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n761), .B2(G326), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1044), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n734), .B1(new_n1037), .B2(new_n1038), .C1(new_n1056), .C2(new_n816), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n685), .A2(new_n802), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1058), .A2(new_n1061), .B1(new_n988), .B2(new_n733), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1030), .A2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n985), .A2(new_n989), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(new_n732), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n959), .A2(new_n802), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n747), .A2(new_n253), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n744), .B1(new_n213), .B2(new_n221), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n734), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(G283), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n264), .B1(new_n782), .B2(new_n1070), .C1(new_n997), .C2(new_n433), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G294), .B2(new_n768), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n772), .A2(new_n783), .B1(new_n618), .B2(new_n778), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT115), .Z(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n1046), .C2(new_n760), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G317), .A2(new_n766), .B1(new_n771), .B2(G311), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n777), .A2(G77), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n830), .A2(new_n258), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G68), .B2(new_n793), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G50), .A2(new_n773), .B1(new_n768), .B2(new_n293), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n823), .C2(new_n760), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G150), .A2(new_n766), .B1(new_n771), .B2(G159), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1075), .A2(new_n1077), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n1085), .B2(new_n740), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1065), .B1(new_n1066), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n988), .A2(new_n728), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1064), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n694), .A3(new_n990), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  AOI211_X1 g0892(.A(new_n922), .B(new_n882), .C1(new_n722), .C2(new_n724), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n931), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n725), .A2(G330), .A3(new_n812), .A4(new_n931), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT116), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n933), .A2(new_n936), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n928), .B1(new_n1099), .B2(new_n931), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n926), .B2(new_n929), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n679), .B(new_n882), .C1(new_n709), .C2(new_n702), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n931), .B1(new_n1102), .B2(new_n935), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n912), .A2(new_n869), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n927), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1098), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1095), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n1098), .C1(new_n1101), .C2(new_n1105), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n727), .B1(new_n477), .B2(new_n478), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n940), .A2(new_n1113), .A3(new_n656), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n932), .B1(new_n726), .B2(new_n882), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1099), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1102), .A2(new_n935), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1118), .A3(new_n1095), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1112), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .A4(new_n1120), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n694), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n734), .B1(new_n298), .B2(new_n840), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n742), .B1(new_n926), .B2(new_n929), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1078), .B1(new_n221), .B2(new_n767), .C1(new_n997), .C2(new_n256), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n761), .B2(G294), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n794), .A2(new_n264), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT118), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n433), .A2(new_n772), .B1(new_n770), .B2(new_n618), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G283), .B2(new_n766), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT119), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n264), .B1(new_n777), .B2(G159), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n997), .B2(new_n202), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n782), .A2(new_n822), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT53), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n767), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1136), .B(new_n1141), .C1(G137), .C2(new_n773), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1137), .A2(new_n1138), .B1(new_n819), .B2(new_n770), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G128), .B2(new_n766), .ZN(new_n1144));
  INV_X1    g0944(.A(G125), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1144), .C1(new_n1145), .C2(new_n760), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1133), .A2(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1134), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1125), .B(new_n1126), .C1(new_n740), .C2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n733), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1124), .A2(KEYINPUT120), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1114), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1123), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n870), .A2(new_n879), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n915), .ZN(new_n1158));
  AND4_X1   g0958(.A1(new_n914), .A2(new_n916), .A3(new_n1104), .A4(new_n893), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n914), .B1(new_n913), .B2(new_n916), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n939), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n908), .A2(new_n917), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1164), .A2(new_n939), .A3(G330), .A4(new_n1158), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n473), .A2(new_n423), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n409), .A2(new_n855), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT121), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  AND2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1163), .A2(new_n1165), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1165), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n939), .B1(new_n918), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1156), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1156), .A2(new_n1178), .A3(KEYINPUT57), .A4(new_n1174), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n694), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1173), .A2(new_n742), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n782), .A2(new_n1140), .B1(new_n822), .B2(new_n778), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G128), .A2(new_n771), .B1(new_n768), .B2(G137), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n819), .B2(new_n772), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G125), .C2(new_n766), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n260), .B(new_n310), .C1(new_n997), .C2(new_n1011), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n761), .B2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n264), .A2(new_n310), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1041), .A2(new_n1009), .A3(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n219), .B2(new_n997), .C1(new_n760), .C2(new_n1070), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n790), .A2(new_n618), .B1(new_n221), .B2(new_n772), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n433), .A2(new_n770), .B1(new_n767), .B2(new_n429), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1195), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1203));
  AND4_X1   g1003(.A1(new_n1194), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n734), .B1(G50), .B2(new_n840), .C1(new_n1204), .C2(new_n816), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1184), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1163), .A2(new_n1165), .A3(new_n1173), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1173), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1206), .B1(new_n1209), .B2(new_n733), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1183), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n733), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n734), .B1(G68), .B2(new_n840), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1008), .B(new_n264), .C1(new_n429), .C2(new_n778), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G97), .B2(new_n793), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G294), .A2(new_n766), .B1(new_n768), .B2(G107), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G116), .A2(new_n773), .B1(new_n771), .B2(G283), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n761), .A2(G303), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n761), .A2(G128), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n258), .B1(new_n782), .B2(new_n1011), .C1(new_n997), .C2(new_n219), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n790), .A2(new_n819), .B1(new_n772), .B2(new_n1140), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT122), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n767), .A2(new_n822), .B1(new_n202), .B2(new_n778), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1002), .A2(G137), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1220), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1214), .B1(new_n1229), .B2(new_n740), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n931), .B2(new_n742), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1213), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1212), .A2(new_n1155), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1121), .A2(new_n972), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(G381));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1091), .A2(new_n844), .A3(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(G381), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1124), .A2(new_n1151), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G387), .A2(new_n1239), .A3(new_n1240), .A4(G375), .ZN(G407));
  NAND3_X1  g1041(.A1(new_n1178), .A2(new_n733), .A3(new_n1174), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1184), .B2(new_n1205), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1028), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1182), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n678), .A2(G213), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  NAND2_X1  g1050(.A1(new_n1234), .A2(KEYINPUT60), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1234), .A2(new_n1253), .A3(KEYINPUT60), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1212), .B2(new_n1155), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n694), .A3(new_n1121), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1260), .B2(new_n1233), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1262), .A2(new_n844), .A3(new_n1232), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1248), .A2(G2897), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(G384), .A3(new_n1233), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n844), .B1(new_n1262), .B2(new_n1232), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(G2897), .A3(new_n1248), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1153), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1124), .A2(new_n1151), .A3(KEYINPUT120), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1183), .A2(new_n1273), .A3(new_n1274), .A4(new_n1210), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1156), .A2(new_n1178), .A3(new_n972), .A4(new_n1174), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1209), .A2(KEYINPUT123), .A3(new_n972), .A4(new_n1156), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1210), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1246), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1275), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1247), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1283), .ZN(new_n1284));
  XOR2_X1   g1084(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1283), .B2(new_n1269), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n992), .A2(new_n1025), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n804), .B1(new_n1030), .B2(new_n1062), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT113), .B1(new_n1237), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1087), .A2(new_n1090), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1237), .A2(new_n1288), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1026), .B(new_n1290), .C1(new_n1091), .C2(new_n1292), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1248), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1284), .A2(new_n1286), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1271), .B2(new_n1298), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1245), .A2(G378), .B1(new_n1280), .B2(new_n1246), .ZN(new_n1303));
  NOR4_X1   g1103(.A1(new_n1303), .A2(KEYINPUT62), .A3(new_n1248), .A4(new_n1269), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1298), .B2(new_n1264), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1302), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1307), .B2(new_n1297), .ZN(G405));
  OAI21_X1  g1108(.A(new_n1275), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT126), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1267), .A2(new_n1311), .A3(new_n1268), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1275), .B(new_n1312), .C1(new_n1240), .C2(new_n1245), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1296), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1296), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AOI211_X1 g1119(.A(KEYINPUT127), .B(new_n1296), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


