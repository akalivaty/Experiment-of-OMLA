//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(G116), .B(G119), .Z(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT2), .B(G113), .Z(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n194), .A3(KEYINPUT71), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n192), .A2(KEYINPUT71), .A3(new_n193), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT64), .A3(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT0), .B(G128), .Z(new_n206));
  AND3_X1   g020(.A1(new_n205), .A2(KEYINPUT65), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n205), .B2(new_n206), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n214), .A2(G137), .B1(KEYINPUT67), .B2(KEYINPUT11), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n214), .A2(G137), .B1(KEYINPUT67), .B2(KEYINPUT11), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n220), .A3(new_n217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n200), .B2(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n203), .A3(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .A4(new_n202), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n226), .A2(new_n229), .A3(G128), .A4(new_n202), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n205), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  OR3_X1    g048(.A1(new_n214), .A2(KEYINPUT69), .A3(G137), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n214), .A2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n212), .B2(G134), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n235), .B(G131), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n221), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n205), .A2(new_n206), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n227), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n216), .A2(new_n220), .A3(new_n217), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n220), .B1(new_n216), .B2(new_n217), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n241), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n209), .A2(new_n222), .A3(KEYINPUT68), .A4(new_n227), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n221), .A2(new_n238), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n221), .B2(new_n238), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n250), .A2(new_n251), .B1(new_n255), .B2(new_n234), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n198), .B(new_n240), .C1(new_n256), .C2(KEYINPUT30), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT31), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n228), .A2(new_n197), .A3(new_n239), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n228), .A2(KEYINPUT72), .A3(new_n197), .A4(new_n239), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(G101), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n265), .B(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n257), .A2(new_n258), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n250), .A2(new_n251), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n255), .A2(new_n234), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT76), .B(new_n198), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n256), .B2(new_n197), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n281), .A3(new_n263), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n272), .A2(new_n273), .B1(new_n284), .B2(new_n269), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n257), .A2(new_n263), .A3(new_n269), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n289), .A3(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT77), .B(new_n188), .C1(new_n285), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n286), .A2(new_n289), .A3(KEYINPUT31), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n286), .B2(KEYINPUT31), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n283), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n275), .ZN(new_n298));
  INV_X1    g112(.A(new_n269), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n270), .B(new_n271), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT77), .B1(new_n302), .B2(new_n188), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n269), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n257), .A2(new_n263), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n276), .A2(KEYINPUT78), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n276), .A2(KEYINPUT78), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n228), .A2(new_n239), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n198), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n263), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n310), .B(new_n311), .C1(new_n314), .C2(new_n274), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n269), .A2(KEYINPUT29), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n308), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT32), .B(new_n188), .C1(new_n285), .C2(new_n291), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT79), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n302), .A2(new_n321), .A3(KEYINPUT32), .A4(new_n188), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n304), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  INV_X1    g139(.A(G128), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(G119), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n328), .A2(KEYINPUT23), .A3(G128), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n327), .A2(new_n329), .B1(G119), .B2(new_n326), .ZN(new_n330));
  XNOR2_X1  g144(.A(G119), .B(G128), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  OAI22_X1  g146(.A1(new_n330), .A2(G110), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n336));
  AND3_X1   g150(.A1(KEYINPUT80), .A2(G125), .A3(G140), .ZN(new_n337));
  AOI21_X1  g151(.A(G140), .B1(KEYINPUT80), .B2(G125), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(KEYINPUT16), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT80), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(KEYINPUT80), .A2(G125), .A3(G140), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n342), .A3(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT81), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n339), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G146), .ZN(new_n349));
  OAI221_X1 g163(.A(KEYINPUT82), .B1(new_n331), .B2(new_n332), .C1(new_n330), .C2(G110), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n203), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n335), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n339), .B(new_n203), .C1(new_n345), .C2(new_n347), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n330), .A2(G110), .B1(new_n331), .B2(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT83), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT22), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(G137), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT84), .Z(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n357), .A3(new_n362), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OR3_X1    g180(.A1(new_n366), .A2(KEYINPUT25), .A3(G902), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(G234), .B2(new_n309), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT25), .B1(new_n366), .B2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(G902), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n365), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G140), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n267), .A2(G227), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G104), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(G107), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n384), .A2(G104), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n381), .A2(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n226), .A2(new_n202), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n232), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n394), .B2(new_n230), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(KEYINPUT85), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(KEYINPUT85), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n380), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n209), .A2(new_n227), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n392), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n234), .A2(new_n405), .A3(KEYINPUT10), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT86), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n404), .A3(new_n409), .A4(new_n406), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n249), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n222), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n379), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n379), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n396), .A2(new_n397), .B1(new_n234), .B2(new_n405), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n415), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT12), .B1(new_n415), .B2(new_n222), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n408), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n222), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n414), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n416), .A2(new_n417), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n379), .B1(new_n425), .B2(new_n412), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n426), .A3(G469), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n420), .A2(new_n309), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n421), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT9), .B(G234), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G221), .B1(new_n432), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n403), .A2(new_n195), .A3(new_n196), .A4(new_n401), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT5), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n328), .A3(G116), .ZN(new_n438));
  OAI211_X1 g252(.A(G113), .B(new_n438), .C1(new_n189), .C2(new_n437), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n405), .A2(new_n194), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT87), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n440), .A3(new_n442), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n447), .A2(new_n441), .A3(new_n448), .A4(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(new_n443), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n436), .B2(new_n440), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n451), .B2(new_n448), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n446), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G125), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n230), .A2(new_n233), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n246), .A2(G125), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n456), .B2(new_n460), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n435), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT88), .B1(new_n444), .B2(KEYINPUT6), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n447), .A3(new_n448), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT90), .A4(new_n446), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n456), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n456), .A2(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n460), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n458), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(new_n460), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n458), .A2(KEYINPUT93), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n479), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n458), .A2(KEYINPUT93), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n439), .A2(new_n194), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n392), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n440), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT91), .B(KEYINPUT8), .Z(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n442), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n481), .A2(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n488), .A3(new_n445), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n472), .A2(new_n309), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n465), .B2(new_n471), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n491), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n266), .A2(new_n267), .A3(G214), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n200), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n349), .A2(new_n501), .A3(new_n354), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n499), .B(G143), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(G131), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n349), .A2(new_n501), .A3(KEYINPUT95), .A4(new_n354), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n381), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n513), .B2(new_n220), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n500), .A2(KEYINPUT18), .A3(G131), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n343), .A2(new_n344), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n352), .B1(new_n516), .B2(new_n203), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT96), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n510), .A2(new_n521), .A3(new_n512), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n505), .B(new_n220), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n506), .A2(KEYINPUT94), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n351), .A2(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(KEYINPUT19), .B2(new_n516), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(G146), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n526), .A2(new_n527), .A3(new_n349), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n518), .ZN(new_n532));
  INV_X1    g346(.A(new_n512), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G475), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n309), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n512), .B1(new_n510), .B2(new_n518), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n520), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g355(.A(G475), .B1(new_n541), .B2(G902), .ZN(new_n542));
  AOI21_X1  g356(.A(G475), .B1(new_n523), .B2(new_n534), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n309), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n200), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n326), .A2(G143), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n214), .ZN(new_n549));
  INV_X1    g363(.A(G116), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT14), .A3(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(G116), .B(G122), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(G107), .B(new_n551), .C1(new_n553), .C2(KEYINPUT14), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n549), .B(new_n554), .C1(G107), .C2(new_n553), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT13), .B1(new_n200), .B2(G128), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n547), .C1(new_n559), .C2(new_n546), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT98), .A3(G134), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n552), .B(new_n384), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n548), .B2(new_n214), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n560), .B2(G134), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n555), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n432), .A2(new_n368), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n555), .B(new_n568), .C1(new_n563), .C2(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT99), .B1(new_n572), .B2(new_n309), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n574), .B(G902), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT15), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(G478), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n572), .B(new_n309), .C1(KEYINPUT15), .C2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(G234), .A2(G237), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(G952), .A3(new_n267), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT21), .B(G898), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(G902), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n545), .A2(new_n581), .A3(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n434), .A2(new_n498), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n324), .A2(new_n375), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  OAI21_X1  g408(.A(new_n188), .B1(new_n285), .B2(new_n291), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n292), .ZN(new_n598));
  INV_X1    g412(.A(new_n433), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n428), .B1(new_n419), .B2(new_n420), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n427), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n302), .A2(new_n309), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n598), .A2(new_n375), .A3(new_n601), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n494), .A2(new_n491), .A3(new_n489), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n491), .B1(new_n494), .B2(new_n489), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n497), .B(new_n590), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n573), .A2(new_n575), .A3(G478), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n560), .A2(G134), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n562), .B(new_n561), .C1(new_n611), .C2(new_n565), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT100), .B1(new_n612), .B2(new_n555), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n572), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n610), .B1(new_n567), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n571), .A3(new_n570), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n579), .A2(G902), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n609), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n608), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n607), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n604), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G6));
  OR2_X1    g440(.A1(new_n581), .A2(new_n608), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n607), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT35), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT102), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n359), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n372), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n371), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n592), .A2(new_n598), .A3(new_n603), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT37), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G110), .ZN(G12));
  NOR2_X1   g453(.A1(new_n434), .A2(new_n498), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n583), .B1(new_n587), .B2(G900), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n324), .A2(new_n640), .A3(new_n636), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  XOR2_X1   g459(.A(new_n641), .B(KEYINPUT39), .Z(new_n646));
  NOR2_X1   g460(.A1(new_n434), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n496), .B(KEYINPUT38), .Z(new_n650));
  INV_X1    g464(.A(new_n314), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n309), .B1(new_n651), .B2(new_n269), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n306), .A2(new_n299), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n304), .A2(new_n323), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n497), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n545), .A2(new_n581), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n649), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n636), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n659), .B(new_n660), .C1(KEYINPUT40), .C2(new_n648), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NOR2_X1   g476(.A1(new_n621), .A2(new_n642), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n324), .A2(new_n640), .A3(new_n636), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  AOI22_X1  g480(.A1(new_n598), .A2(new_n187), .B1(new_n320), .B2(new_n322), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n374), .B1(new_n667), .B2(new_n318), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n419), .A2(new_n420), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n421), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n599), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n622), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n324), .A2(new_n375), .A3(new_n622), .A4(new_n671), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT41), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G113), .ZN(G15));
  NAND4_X1  g492(.A1(new_n324), .A2(new_n375), .A3(new_n628), .A4(new_n671), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  INV_X1    g494(.A(new_n591), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n670), .A2(new_n498), .A3(new_n599), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n324), .A2(new_n681), .A3(new_n636), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT105), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NAND2_X1  g499(.A1(new_n315), .A2(new_n299), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n301), .A2(new_n287), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n188), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n603), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n375), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(KEYINPUT106), .A3(new_n375), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n657), .A2(new_n496), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n590), .A3(new_n671), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NAND3_X1  g512(.A1(new_n603), .A2(new_n636), .A3(new_n688), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n663), .A3(new_n682), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT107), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n454), .ZN(G27));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n427), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT108), .A4(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n600), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n433), .A2(new_n497), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n496), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n324), .A2(new_n375), .A3(new_n663), .A4(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n595), .A2(new_n187), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n318), .A3(new_n319), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n375), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n663), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n709), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT109), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n721), .B(new_n718), .C1(new_n711), .C2(new_n712), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n220), .ZN(G33));
  NAND4_X1  g538(.A1(new_n668), .A2(KEYINPUT110), .A3(new_n643), .A4(new_n710), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n324), .A2(new_n375), .A3(new_n643), .A4(new_n710), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  NAND2_X1  g544(.A1(new_n424), .A2(new_n426), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n429), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n421), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT111), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT111), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n428), .B1(new_n732), .B2(G469), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n736), .B(new_n737), .C1(KEYINPUT46), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n433), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n646), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n545), .A2(new_n620), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT43), .Z(new_n743));
  AOI21_X1  g557(.A(new_n660), .B1(new_n598), .B2(new_n603), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n656), .B(new_n496), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n741), .B(new_n747), .C1(new_n746), .C2(new_n745), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n740), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n433), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n324), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n496), .A2(new_n656), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n374), .A3(new_n663), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n607), .B2(new_n621), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n609), .A2(new_n619), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT20), .B1(new_n543), .B2(new_n309), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n520), .A2(new_n522), .B1(new_n533), .B2(new_n532), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n761), .A2(new_n538), .A3(G475), .A4(G902), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n763), .B2(new_n542), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n656), .B1(new_n493), .B2(new_n495), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n590), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n604), .A2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n593), .A2(new_n769), .A3(KEYINPUT113), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT113), .B1(new_n593), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n637), .A2(new_n629), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n581), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n608), .A2(new_n774), .A3(new_n642), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n324), .A2(new_n601), .A3(new_n754), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n710), .A2(new_n689), .A3(new_n663), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n728), .A2(new_n725), .B1(new_n778), .B2(new_n636), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n433), .A2(new_n707), .A3(new_n660), .A4(new_n496), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n655), .A2(new_n780), .A3(new_n641), .A4(new_n657), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n644), .A2(new_n781), .A3(new_n664), .A4(new_n701), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n660), .B1(new_n667), .B2(new_n318), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n640), .A2(new_n643), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n682), .A2(new_n663), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(new_n700), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n664), .A4(new_n781), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n773), .A2(new_n779), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n672), .A2(new_n675), .B1(new_n694), .B2(new_n696), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n679), .A2(new_n683), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n791), .B(new_n792), .C1(new_n720), .C2(new_n722), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n757), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n673), .A2(new_n674), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n673), .A2(new_n674), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n792), .B(new_n697), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n718), .B1(new_n711), .B2(new_n712), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n757), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n593), .A2(new_n769), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n593), .A2(new_n769), .A3(KEYINPUT113), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n629), .A3(new_n637), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n778), .A2(new_n636), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n729), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n789), .A2(new_n783), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n794), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n723), .A2(new_n797), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n807), .A4(new_n808), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n813), .B2(new_n794), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n794), .A2(new_n809), .A3(new_n810), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT115), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n814), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(KEYINPUT114), .A3(new_n817), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  INV_X1    g636(.A(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n751), .A2(new_n752), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n751), .A2(KEYINPUT116), .A3(new_n752), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n669), .A2(new_n599), .A3(new_n421), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n694), .A2(new_n584), .A3(new_n743), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n754), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n834));
  INV_X1    g648(.A(new_n655), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n375), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n671), .A2(new_n584), .A3(new_n754), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n837), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n835), .A3(KEYINPUT118), .A4(new_n375), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n545), .A3(new_n759), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(KEYINPUT119), .A3(new_n545), .A4(new_n759), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n650), .A2(new_n671), .A3(new_n656), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT117), .Z(new_n848));
  NAND2_X1  g662(.A1(new_n831), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n831), .A2(new_n848), .A3(KEYINPUT50), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n839), .A2(new_n743), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n851), .A2(new_n852), .B1(new_n700), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n846), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT51), .B1(new_n833), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n751), .A2(new_n752), .A3(new_n829), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n832), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n846), .A2(new_n859), .A3(KEYINPUT51), .A4(new_n855), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n831), .A2(new_n682), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n853), .A2(new_n716), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT48), .Z(new_n863));
  INV_X1    g677(.A(G952), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n864), .B(G953), .C1(new_n841), .C2(new_n764), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n861), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n819), .A2(new_n824), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n267), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n819), .A2(new_n824), .A3(KEYINPUT120), .A4(new_n867), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n708), .B1(new_n670), .B2(KEYINPUT49), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n375), .B1(new_n670), .B2(KEYINPUT49), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n742), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n835), .A2(new_n650), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n877), .ZN(G75));
  AOI21_X1  g692(.A(new_n309), .B1(new_n794), .B2(new_n809), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n453), .B(new_n470), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n880), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n267), .A2(G952), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(G51));
  AOI21_X1  g699(.A(new_n810), .B1(new_n794), .B2(new_n809), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n811), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n428), .B(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n413), .A2(new_n418), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n879), .A2(G469), .A3(new_n732), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n884), .B1(new_n893), .B2(new_n894), .ZN(G54));
  AND3_X1   g709(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n535), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT122), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n535), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n898), .A2(new_n884), .A3(new_n899), .ZN(G60));
  XNOR2_X1  g714(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n887), .A2(new_n614), .A3(new_n617), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n819), .A2(new_n824), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n614), .A2(new_n617), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n884), .B(new_n905), .C1(new_n907), .C2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n794), .B2(new_n809), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n884), .B1(new_n912), .B2(new_n634), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n366), .B(KEYINPUT124), .Z(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n586), .B2(new_n457), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n797), .A2(new_n804), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n453), .B1(G898), .B2(new_n267), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(new_n755), .A2(new_n748), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n723), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n741), .A2(new_n375), .A3(new_n695), .A4(new_n715), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n644), .A2(new_n664), .A3(new_n701), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n924), .A2(new_n729), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n267), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n240), .B1(new_n256), .B2(KEYINPUT30), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT125), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n529), .ZN(new_n931));
  NAND2_X1  g745(.A1(G900), .A2(G953), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n926), .A2(new_n661), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT62), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n627), .A2(new_n621), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n668), .A2(new_n647), .A3(new_n754), .A4(new_n936), .ZN(new_n937));
  AND4_X1   g751(.A1(new_n748), .A2(new_n935), .A3(new_n755), .A4(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n939), .B2(new_n931), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G72));
  INV_X1    g756(.A(new_n653), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n918), .ZN(new_n944));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n307), .B(KEYINPUT127), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n923), .A2(new_n918), .A3(new_n927), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n813), .A2(new_n794), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n307), .A2(new_n951), .A3(new_n943), .A4(new_n946), .ZN(new_n952));
  NOR4_X1   g766(.A1(new_n947), .A2(new_n884), .A3(new_n950), .A4(new_n952), .ZN(G57));
endmodule


