//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT71), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n203), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT24), .B1(new_n215), .B2(KEYINPUT65), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n210), .B1(new_n217), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT23), .B2(new_n218), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(KEYINPUT25), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n214), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n237), .A3(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G176gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT23), .A4(new_n220), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n215), .A2(new_n232), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  INV_X1    g043(.A(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n246), .A3(new_n211), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n247), .A3(new_n223), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n238), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n215), .B1(new_n222), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n218), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT27), .B(G183gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n245), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n259), .A4(new_n245), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n251), .A2(new_n252), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n251), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n209), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n252), .A3(new_n264), .ZN(new_n271));
  INV_X1    g070(.A(new_n209), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n256), .A2(new_n262), .A3(new_n263), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n230), .A2(new_n237), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n274), .A2(new_n210), .B1(new_n249), .B2(new_n248), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(new_n238), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n271), .B(new_n272), .C1(new_n276), .C2(new_n266), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT72), .B(new_n209), .C1(new_n265), .C2(new_n267), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT73), .ZN(new_n281));
  XNOR2_X1  g080(.A(G64gat), .B(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT74), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n270), .A2(new_n277), .A3(new_n278), .A4(new_n283), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G1gat), .B(G29gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT0), .ZN(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n296), .A2(G155gat), .A3(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT76), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n295), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(KEYINPUT2), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n301), .A2(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n295), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT76), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n296), .B1(G155gat), .B2(G162gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT2), .B1(new_n317), .B2(new_n298), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n306), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n299), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n295), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n305), .A2(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n309), .A2(new_n314), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n327), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(G127gat), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n329), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n327), .B2(KEYINPUT1), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  INV_X1    g139(.A(G134gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n332), .A2(G120gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n330), .A2(G113gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n335), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT4), .B1(new_n326), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n340), .B1(new_n339), .B2(new_n344), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(KEYINPUT78), .A2(new_n323), .B1(new_n321), .B2(new_n295), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n318), .A2(new_n320), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n307), .A2(new_n308), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n313), .B2(KEYINPUT77), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n358), .A3(new_n346), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n347), .B1(new_n360), .B2(KEYINPUT4), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n301), .A2(new_n302), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n314), .A3(new_n354), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n352), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n350), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n294), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n369), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n373), .B(new_n374), .C1(new_n326), .C2(new_n346), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n364), .B(new_n352), .C1(new_n348), .C2(new_n349), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT81), .B1(new_n376), .B2(KEYINPUT4), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n374), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n350), .A2(new_n356), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n359), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n369), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n371), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  INV_X1    g186(.A(new_n372), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT4), .B1(new_n350), .B2(new_n356), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n373), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n376), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT4), .B1(new_n357), .B2(new_n359), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n368), .B1(new_n382), .B2(new_n383), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n395), .B1(new_n361), .B2(new_n370), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n386), .B(new_n387), .C1(new_n396), .C2(new_n293), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n361), .A2(new_n370), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n380), .B2(new_n385), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n294), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n289), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n271), .B1(new_n276), .B2(new_n266), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT72), .B1(new_n402), .B2(new_n209), .ZN(new_n403));
  INV_X1    g202(.A(new_n278), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n277), .A4(new_n283), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n288), .A2(KEYINPUT75), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n287), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n401), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n420), .B2(new_n416), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n366), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n209), .B1(new_n423), .B2(KEYINPUT29), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n424), .A2(G228gat), .A3(G233gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n209), .A2(KEYINPUT29), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n356), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n362), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT84), .B(new_n356), .C1(new_n426), .C2(KEYINPUT3), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT85), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n425), .A2(new_n433), .A3(new_n429), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n208), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n436), .A2(new_n202), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n436), .B2(new_n202), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n365), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n356), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n424), .A2(new_n441), .B1(G228gat), .B2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n422), .B1(new_n435), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n442), .B(new_n421), .C1(new_n432), .C2(new_n434), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n251), .A2(new_n264), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(new_n350), .ZN(new_n448));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT33), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT34), .B1(new_n448), .B2(new_n450), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n447), .B(new_n346), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT34), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n450), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n458), .B(new_n461), .C1(new_n451), .C2(new_n456), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n463), .B2(new_n467), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n411), .A2(new_n413), .A3(new_n446), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n288), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n473), .A2(KEYINPUT30), .B1(new_n279), .B2(new_n285), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n409), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n293), .B(KEYINPUT87), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n386), .B(new_n387), .C1(new_n396), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n400), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT90), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n471), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n444), .A2(new_n445), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT35), .ZN(new_n488));
  AOI22_X1  g287(.A1(KEYINPUT35), .A2(new_n472), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n397), .A2(new_n400), .ZN(new_n490));
  AND4_X1   g289(.A1(new_n412), .A2(new_n490), .A3(new_n409), .A4(new_n474), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n412), .B1(new_n401), .B2(new_n409), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n357), .A2(new_n359), .A3(new_n369), .A4(new_n381), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(KEYINPUT39), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n374), .B1(new_n357), .B2(new_n359), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n362), .A2(new_n350), .A3(new_n366), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n496), .A2(new_n347), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n498), .B2(new_n369), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g299(.A(new_n347), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n367), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n383), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n504), .A3(new_n478), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n499), .A2(new_n504), .A3(KEYINPUT40), .A4(new_n478), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n399), .A2(new_n477), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n475), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n268), .A2(new_n277), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n265), .A2(new_n267), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n272), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(KEYINPUT37), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT37), .B1(new_n514), .B2(new_n272), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n270), .A3(new_n278), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n284), .A2(KEYINPUT38), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n407), .A2(new_n520), .A3(new_n408), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n279), .A2(KEYINPUT37), .ZN(new_n522));
  INV_X1    g321(.A(new_n283), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT38), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n400), .A3(new_n479), .A4(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n526), .A3(new_n446), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT89), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n469), .B2(new_n470), .ZN(new_n530));
  INV_X1    g329(.A(new_n470), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(KEYINPUT36), .A3(new_n468), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n511), .A2(new_n526), .A3(new_n534), .A4(new_n446), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n489), .B1(new_n493), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT12), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT14), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT14), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT92), .Z(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT93), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT15), .B(new_n552), .C1(new_n550), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT17), .ZN(new_n562));
  XOR2_X1   g361(.A(G15gat), .B(G22gat), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G1gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565));
  INV_X1    g364(.A(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT16), .ZN(new_n567));
  OAI221_X1 g366(.A(new_n564), .B1(new_n565), .B2(G8gat), .C1(new_n563), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(G8gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n561), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(KEYINPUT18), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n544), .B1(new_n576), .B2(KEYINPUT95), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(KEYINPUT18), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n570), .B(new_n573), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n572), .B(KEYINPUT13), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n537), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT98), .B(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n589), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n594), .A2(KEYINPUT99), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT8), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n594), .B2(KEYINPUT99), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n595), .A2(new_n597), .B1(new_n590), .B2(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n602), .A3(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n588), .B1(new_n573), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n562), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G57gat), .B(G64gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G71gat), .B(G78gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n570), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n298), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n624), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G127gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n627), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  INV_X1    g439(.A(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n604), .B(new_n622), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(KEYINPUT10), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n604), .A2(new_n622), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT10), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n642), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n639), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n639), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n652), .B2(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n636), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n587), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n490), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g460(.A1(new_n537), .A2(new_n476), .A3(new_n586), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n657), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT103), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  MUX2_X1   g465(.A(KEYINPUT103), .B(new_n665), .S(new_n666), .Z(new_n667));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n663), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n669), .B2(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(G8gat), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n673), .A3(new_n471), .ZN(new_n674));
  INV_X1    g473(.A(new_n533), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n658), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n676), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n487), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n678), .B(new_n679), .ZN(new_n684));
  INV_X1    g483(.A(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(G1327gat));
  NAND2_X1  g486(.A1(new_n536), .A2(new_n493), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n485), .A2(new_n488), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n656), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n634), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n586), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n692), .A2(new_n614), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n545), .A3(new_n659), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n493), .A2(KEYINPUT106), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n535), .A2(new_n533), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n701), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n699), .A2(new_n528), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n691), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n691), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n615), .A2(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n537), .B2(new_n615), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n695), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n712), .B2(new_n490), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G29gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n490), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n698), .B1(new_n714), .B2(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n476), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n694), .A2(new_n615), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n662), .A2(new_n546), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n717), .B(new_n722), .C1(new_n720), .C2(new_n719), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n724), .A3(new_n471), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n712), .A2(new_n533), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT47), .B(new_n725), .C1(new_n726), .C2(new_n724), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n446), .B2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n487), .A2(KEYINPUT110), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n587), .A2(new_n718), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n712), .A2(new_n446), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n734), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT48), .B(new_n736), .C1(new_n737), .C2(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NOR3_X1   g541(.A1(new_n636), .A2(new_n693), .A3(new_n585), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n705), .A2(new_n707), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n490), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(G57gat), .Z(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(KEYINPUT111), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n705), .A2(new_n748), .A3(new_n707), .A4(new_n743), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n475), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n747), .A2(new_n675), .A3(new_n749), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n744), .A2(G71gat), .A3(new_n486), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1334gat));
  NAND3_X1  g558(.A1(new_n747), .A2(new_n487), .A3(new_n749), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g560(.A(KEYINPUT113), .B1(new_n585), .B2(new_n635), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n583), .A2(new_n634), .A3(new_n763), .A4(new_n584), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n656), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n711), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n490), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n411), .A2(new_n413), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n701), .B1(new_n771), .B2(new_n487), .ZN(new_n772));
  INV_X1    g571(.A(new_n702), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n489), .B1(new_n774), .B2(new_n536), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n765), .A2(new_n614), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n704), .A3(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n656), .A2(new_n590), .A3(new_n659), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n769), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n768), .B2(new_n476), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n785), .A3(new_n779), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT114), .B(new_n770), .C1(new_n775), .C2(new_n776), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n693), .A2(G92gat), .A3(new_n476), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(new_n780), .B2(new_n788), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n768), .B2(new_n533), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n693), .A2(G99gat), .A3(new_n486), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT116), .Z(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n781), .B2(new_n800), .ZN(G1338gat));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n703), .A2(new_n706), .A3(new_n691), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n706), .B1(new_n703), .B2(new_n691), .ZN(new_n805));
  INV_X1    g604(.A(new_n708), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n692), .B2(new_n614), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n487), .B(new_n767), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n693), .A2(G106gat), .A3(new_n446), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT117), .Z(new_n813));
  NAND3_X1  g612(.A1(new_n786), .A2(new_n787), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n803), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n766), .B1(new_n709), .B2(new_n710), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n487), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n780), .A2(new_n812), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n803), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n802), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n786), .A2(new_n787), .A3(new_n813), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT53), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n811), .A2(new_n803), .A3(new_n819), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT118), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n644), .A2(new_n642), .A3(new_n646), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n648), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n639), .B1(new_n647), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n834), .A2(new_n655), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n585), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n582), .A2(new_n543), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n579), .A2(new_n580), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n838), .B1(new_n542), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n656), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n614), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n842), .A2(new_n836), .A3(new_n614), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n634), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n657), .A2(new_n586), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n487), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n471), .A2(new_n659), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n475), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n585), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n332), .A2(KEYINPUT119), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n332), .A2(KEYINPUT119), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n851), .B2(new_n852), .ZN(G1340gat));
  NAND2_X1  g654(.A1(new_n848), .A2(new_n850), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n693), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(new_n330), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n635), .A3(new_n850), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT120), .ZN(new_n860));
  XOR2_X1   g659(.A(KEYINPUT68), .B(G127gat), .Z(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1342gat));
  NOR3_X1   g661(.A1(new_n615), .A2(new_n475), .A3(new_n849), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(KEYINPUT56), .A3(new_n341), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n864), .B2(new_n341), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n865), .A2(new_n866), .B1(new_n341), .B2(new_n864), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n675), .A2(new_n490), .A3(new_n475), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n586), .A2(new_n305), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n487), .A2(KEYINPUT57), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n846), .A2(KEYINPUT122), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n846), .A2(KEYINPUT122), .B1(new_n586), .B2(new_n657), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n446), .B1(new_n846), .B2(new_n847), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n868), .B(new_n869), .C1(new_n873), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n585), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n305), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT123), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n882), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT123), .B(new_n884), .C1(new_n878), .C2(new_n880), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(new_n874), .ZN(new_n887));
  INV_X1    g686(.A(new_n868), .ZN(new_n888));
  NOR4_X1   g687(.A1(new_n887), .A2(G148gat), .A3(new_n693), .A4(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT125), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n873), .A2(new_n877), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n888), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n656), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n656), .B1(new_n868), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n896), .B2(new_n868), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n887), .A2(new_n875), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n891), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n890), .B1(new_n895), .B2(new_n902), .ZN(G1345gat));
  AOI21_X1  g702(.A(new_n298), .B1(new_n894), .B2(new_n635), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n887), .A2(G155gat), .A3(new_n634), .A4(new_n888), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  NAND4_X1  g705(.A1(new_n874), .A2(new_n317), .A3(new_n614), .A4(new_n868), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n894), .A2(new_n614), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n909), .B2(new_n317), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n846), .A2(new_n847), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n475), .A2(new_n490), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n486), .A2(new_n487), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n586), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(new_n220), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n656), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G176gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n239), .A2(new_n241), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(G1349gat));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n635), .A3(new_n913), .ZN(new_n921));
  MUX2_X1   g720(.A(new_n257), .B(G183gat), .S(new_n921), .Z(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT60), .ZN(G1350gat));
  OAI22_X1  g722(.A1(new_n914), .A2(new_n615), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n675), .A2(new_n912), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n874), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n874), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n585), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n927), .B1(new_n899), .B2(new_n900), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n585), .A2(G197gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n928), .A2(G204gat), .A3(new_n693), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT62), .ZN(new_n940));
  OAI21_X1  g739(.A(G204gat), .B1(new_n935), .B2(new_n693), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1353gat));
  OAI211_X1 g741(.A(new_n635), .B(new_n927), .C1(new_n899), .C2(new_n900), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n635), .A2(new_n205), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n944), .A2(new_n945), .B1(new_n932), .B2(new_n946), .ZN(G1354gat));
  NAND3_X1  g746(.A1(new_n933), .A2(new_n206), .A3(new_n614), .ZN(new_n948));
  OAI21_X1  g747(.A(G218gat), .B1(new_n935), .B2(new_n615), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1355gat));
endmodule


