//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(new_n213), .B2(new_n212), .ZN(new_n218));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT2), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G155gat), .B(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n224), .A3(new_n222), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n218), .B1(KEYINPUT29), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(KEYINPUT78), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n231), .A2(KEYINPUT78), .B1(G228gat), .B2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n217), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n212), .A2(new_n213), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n216), .A2(KEYINPUT77), .A3(new_n217), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n228), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT72), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n232), .B(new_n233), .C1(new_n241), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(new_n237), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(new_n246), .B2(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(new_n242), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n231), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(G228gat), .A3(G233gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n245), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n206), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n205), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT23), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT24), .ZN(new_n265));
  INV_X1    g064(.A(G169gat), .ZN(new_n266));
  INV_X1    g065(.A(G176gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .A3(new_n264), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  INV_X1    g074(.A(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n268), .A2(KEYINPUT26), .A3(new_n261), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n261), .A2(KEYINPUT26), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n264), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n285), .A2(new_n240), .B1(G226gat), .B2(G233gat), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n272), .A2(new_n273), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n273), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(new_n288), .B1(new_n279), .B2(new_n283), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n218), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n289), .B2(KEYINPUT29), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n246), .C1(new_n290), .C2(new_n289), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT70), .A4(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n305), .A3(new_n301), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n294), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n309), .A2(new_n297), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n298), .A2(new_n301), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313));
  XOR2_X1   g112(.A(G1gat), .B(G29gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT0), .ZN(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT79), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT39), .ZN(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT4), .B1(new_n332), .B2(new_n244), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(new_n226), .A3(new_n329), .A4(new_n228), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n330), .A3(new_n229), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n320), .B(new_n322), .C1(new_n333), .C2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n333), .A2(new_n339), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(new_n321), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n242), .A2(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n334), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n322), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n320), .B1(new_n345), .B2(KEYINPUT80), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(KEYINPUT80), .B2(new_n345), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n319), .B(new_n340), .C1(new_n342), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT40), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n313), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n342), .A2(new_n347), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n319), .A2(new_n340), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(KEYINPUT81), .A3(KEYINPUT40), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n322), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n332), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n322), .B1(new_n334), .B2(new_n335), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n338), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT73), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n356), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR4_X1   g163(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT5), .A4(new_n322), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n318), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n366), .A2(KEYINPUT40), .B1(new_n351), .B2(new_n352), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n354), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n260), .B1(new_n312), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT82), .B1(new_n308), .B2(KEYINPUT37), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT37), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n292), .A2(new_n294), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n297), .B1(new_n308), .B2(KEYINPUT37), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT38), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(KEYINPUT38), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n365), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n317), .ZN(new_n384));
  INV_X1    g183(.A(new_n317), .ZN(new_n385));
  NOR4_X1   g184(.A1(new_n364), .A2(KEYINPUT74), .A3(new_n385), .A4(new_n365), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n381), .B(new_n366), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(KEYINPUT6), .B(new_n385), .C1(new_n364), .C2(new_n365), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT75), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n300), .A2(new_n302), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(new_n387), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n369), .A2(new_n391), .A3(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n332), .A2(new_n285), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n330), .B(KEYINPUT65), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n289), .ZN(new_n398));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT64), .Z(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT68), .ZN(new_n403));
  XOR2_X1   g202(.A(G71gat), .B(G99gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT33), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(KEYINPUT32), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n401), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n401), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n401), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n407), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n398), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n399), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT34), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n407), .C1(new_n412), .C2(new_n417), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT36), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT36), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n310), .A2(new_n311), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n304), .B2(new_n306), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n381), .B1(new_n383), .B2(new_n317), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n383), .A2(new_n317), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT74), .ZN(new_n437));
  INV_X1    g236(.A(new_n386), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n388), .B(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n434), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n432), .B1(new_n442), .B2(new_n260), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n394), .A2(new_n395), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n366), .A2(new_n381), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n437), .B2(new_n438), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n445), .B(new_n434), .C1(new_n447), .C2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n260), .A2(new_n428), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n384), .A2(new_n386), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n389), .B1(new_n452), .B2(new_n435), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n453), .A3(new_n434), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n458));
  NAND2_X1  g257(.A1(G229gat), .A2(G233gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n459), .B(KEYINPUT89), .Z(new_n460));
  AND2_X1   g259(.A1(G43gat), .A2(G50gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(G43gat), .A2(G50gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT85), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G43gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n203), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g265(.A1(G43gat), .A2(G50gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n468), .A3(KEYINPUT15), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n461), .A2(new_n462), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT86), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G36gat), .ZN(new_n474));
  AND2_X1   g273(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n471), .A3(new_n467), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n469), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G22gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G15gat), .ZN(new_n489));
  INV_X1    g288(.A(G15gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G22gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT87), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G8gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT87), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  AOI21_X1  g297(.A(G1gat), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n493), .A3(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT90), .B1(new_n487), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n499), .A2(new_n493), .A3(new_n496), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n499), .B1(new_n493), .B2(new_n496), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n473), .A2(new_n480), .B1(new_n485), .B2(new_n469), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n460), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n465), .A2(new_n467), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n471), .B1(new_n514), .B2(KEYINPUT85), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n468), .A2(new_n515), .B1(new_n480), .B2(new_n484), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n478), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT14), .B(G29gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n474), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n469), .B2(new_n472), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n513), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n481), .A2(KEYINPUT17), .A3(new_n486), .ZN(new_n522));
  AOI211_X1 g321(.A(new_n512), .B(new_n507), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT88), .B1(new_n524), .B2(new_n503), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT18), .B(new_n511), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n487), .A2(new_n503), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n487), .A2(new_n503), .A3(KEYINPUT90), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n509), .B1(new_n507), .B2(new_n508), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n460), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n460), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n528), .B2(new_n529), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n516), .A2(new_n520), .A3(new_n513), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT17), .B1(new_n481), .B2(new_n486), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n503), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n512), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT88), .A3(new_n503), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n526), .B(new_n533), .C1(new_n541), .C2(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT84), .B(G197gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT11), .B(G169gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT12), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT12), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n530), .A2(new_n532), .B1(new_n552), .B2(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n526), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n540), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT18), .B1(new_n557), .B2(new_n511), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n511), .B1(new_n523), .B2(new_n525), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(KEYINPUT92), .A3(new_n526), .A4(new_n555), .ZN(new_n563));
  AOI221_X4 g362(.A(new_n458), .B1(new_n542), .B2(new_n553), .C1(new_n559), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n542), .A2(new_n553), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT93), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n457), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G57gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT94), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n572), .A2(new_n574), .B1(new_n577), .B2(new_n576), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n583), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n583), .A2(KEYINPUT95), .A3(new_n580), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT95), .B1(new_n583), .B2(new_n580), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n582), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n507), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G127gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(G127gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(new_n590), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n220), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n598), .A2(new_n601), .A3(new_n606), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G99gat), .ZN(new_n615));
  INV_X1    g414(.A(G106gat), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT8), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G85gat), .A2(G92gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT97), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT7), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n624), .A3(KEYINPUT7), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n618), .A2(new_n620), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n617), .A3(new_n614), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n619), .B1(new_n629), .B2(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n524), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n633), .A2(new_n508), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G134gat), .B(G162gat), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n637), .B(KEYINPUT99), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI221_X1 g443(.A(new_n639), .B1(KEYINPUT100), .B2(new_n642), .C1(new_n636), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n588), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n579), .B2(new_n581), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n583), .A2(KEYINPUT95), .A3(new_n580), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n579), .A2(KEYINPUT94), .A3(new_n581), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n584), .B1(new_n583), .B2(new_n580), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n658), .A2(new_n628), .A3(new_n630), .A4(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n653), .B1(new_n654), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT102), .Z(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n633), .A2(new_n589), .A3(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n653), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n676));
  INV_X1    g475(.A(new_n653), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n666), .B2(new_n667), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n673), .A3(new_n676), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n610), .A2(new_n652), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n570), .A2(new_n453), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n434), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT104), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n457), .A2(new_n569), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n693));
  INV_X1    g492(.A(new_n687), .ZN(new_n694));
  OAI21_X1  g493(.A(G8gat), .B1(new_n570), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n693), .A2(new_n699), .A3(new_n695), .A4(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(new_n432), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n570), .A2(new_n702), .A3(new_n684), .ZN(new_n703));
  INV_X1    g502(.A(new_n684), .ZN(new_n704));
  INV_X1    g503(.A(new_n428), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n490), .A3(new_n705), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n703), .A2(new_n490), .B1(new_n570), .B2(new_n706), .ZN(G1326gat));
  INV_X1    g506(.A(new_n260), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n570), .A2(new_n708), .A3(new_n684), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n450), .A2(new_n449), .B1(new_n454), .B2(KEYINPUT35), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n442), .A2(new_n260), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n702), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT83), .B1(new_n369), .B2(new_n391), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(new_n395), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n718), .B2(new_n652), .ZN(new_n719));
  INV_X1    g518(.A(new_n453), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n457), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n610), .B(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n565), .A2(new_n566), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n722), .A2(new_n724), .A3(new_n682), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G29gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n610), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n651), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n682), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n453), .A2(G29gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n457), .A2(new_n569), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n727), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n570), .A2(new_n682), .A3(new_n729), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n434), .A2(G36gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n745), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n457), .B2(new_n651), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n712), .B(new_n652), .C1(new_n444), .C2(new_n456), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n312), .A3(new_n725), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G36gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n746), .A2(new_n748), .A3(new_n753), .ZN(G1329gat));
  NAND4_X1  g553(.A1(new_n719), .A2(new_n432), .A3(new_n721), .A4(new_n725), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n464), .A3(new_n705), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1330gat));
  NAND4_X1  g562(.A1(new_n719), .A2(new_n260), .A3(new_n721), .A4(new_n725), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G50gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n740), .A2(new_n203), .A3(new_n260), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT48), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  NOR4_X1   g570(.A1(new_n728), .A2(new_n723), .A3(new_n651), .A4(new_n683), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n457), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n453), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT110), .B(G57gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1332gat));
  INV_X1    g575(.A(new_n773), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n434), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1333gat));
  OR3_X1    g584(.A1(new_n773), .A2(G71gat), .A3(new_n428), .ZN(new_n786));
  OAI21_X1  g585(.A(G71gat), .B1(new_n773), .B2(new_n702), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g588(.A1(new_n777), .A2(new_n260), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g590(.A(new_n652), .B1(new_n444), .B2(new_n456), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n610), .A2(new_n723), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT51), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT112), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT112), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n453), .A2(G85gat), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n796), .A2(new_n682), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n610), .A2(new_n723), .A3(new_n683), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n751), .A2(new_n720), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n612), .B2(new_n801), .ZN(G1336gat));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n719), .A2(new_n312), .A3(new_n721), .A4(new_n800), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n611), .A2(new_n613), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n434), .A2(G92gat), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n682), .B(new_n810), .C1(new_n794), .C2(new_n795), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n803), .A2(new_n804), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n805), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n806), .B2(new_n808), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n805), .B1(new_n815), .B2(new_n811), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n814), .A2(new_n816), .ZN(G1337gat));
  NOR2_X1   g616(.A1(new_n428), .A2(G99gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n796), .A2(new_n682), .A3(new_n797), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n751), .A2(new_n432), .A3(new_n800), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n615), .B2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n719), .A2(new_n260), .A3(new_n721), .A4(new_n800), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n708), .A2(G106gat), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n682), .B(new_n824), .C1(new_n794), .C2(new_n795), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n751), .A2(new_n828), .A3(new_n260), .A4(new_n800), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n829), .A2(new_n830), .A3(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n831), .B2(new_n833), .ZN(G1339gat));
  NOR2_X1   g633(.A1(new_n684), .A2(new_n723), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n666), .A2(new_n667), .A3(new_n677), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n676), .A2(new_n838), .A3(new_n680), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT54), .B(new_n677), .C1(new_n666), .C2(new_n667), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(new_n673), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n678), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT115), .B1(new_n844), .B2(new_n674), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n839), .B(KEYINPUT55), .C1(new_n842), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n681), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n681), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n839), .B1(new_n842), .B2(new_n845), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n504), .A2(new_n510), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n534), .B1(new_n557), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n530), .A2(new_n532), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n550), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n651), .A2(new_n565), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n682), .A2(new_n565), .A3(new_n858), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n854), .B2(new_n724), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n862), .B2(new_n652), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n836), .B1(new_n863), .B2(new_n722), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n450), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n453), .A2(new_n312), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n568), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT117), .Z(new_n869));
  XNOR2_X1  g668(.A(new_n867), .B(KEYINPUT118), .ZN(new_n870));
  INV_X1    g669(.A(G113gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n723), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(G1340gat));
  OAI21_X1  g672(.A(G120gat), .B1(new_n867), .B2(new_n683), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(G120gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n870), .A2(new_n876), .A3(new_n682), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n722), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n867), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n867), .A2(KEYINPUT120), .A3(new_n728), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(G127gat), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT120), .B1(new_n867), .B2(new_n728), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1342gat));
  AOI211_X1 g684(.A(new_n652), .B(new_n867), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n864), .A2(new_n260), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n702), .A2(new_n866), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(G141gat), .A3(new_n568), .ZN(new_n893));
  INV_X1    g692(.A(new_n890), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n864), .B2(new_n260), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n708), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n853), .A2(new_n681), .A3(new_n846), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n723), .A2(new_n458), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n565), .A2(KEYINPUT93), .A3(new_n566), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n861), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n652), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n854), .A2(new_n859), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n610), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n836), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n841), .B1(new_n840), .B2(new_n673), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n844), .A2(KEYINPUT115), .A3(new_n674), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT55), .B1(new_n911), .B2(new_n839), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n847), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n564), .B2(new_n567), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n651), .B1(new_n914), .B2(new_n861), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n907), .B(new_n728), .C1(new_n915), .C2(new_n860), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n898), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n896), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n898), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n728), .B1(new_n915), .B2(new_n860), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n835), .B1(new_n922), .B2(KEYINPUT121), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n916), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n723), .B(new_n894), .C1(new_n920), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n893), .B1(new_n926), .B2(G141gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n929));
  INV_X1    g728(.A(G141gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n895), .B1(new_n924), .B2(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n918), .A2(new_n919), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n890), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n569), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n927), .A2(new_n928), .B1(new_n929), .B2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(G148gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n891), .A2(new_n936), .A3(new_n682), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT59), .B(new_n936), .C1(new_n933), .C2(new_n682), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n569), .A2(new_n684), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n260), .B1(new_n906), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n897), .ZN(new_n943));
  INV_X1    g742(.A(new_n940), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n708), .B1(new_n922), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT124), .B1(new_n945), .B2(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n864), .A2(new_n898), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n682), .A3(new_n894), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n939), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n937), .B1(new_n938), .B2(new_n950), .ZN(G1345gat));
  NAND3_X1  g750(.A1(new_n891), .A2(new_n220), .A3(new_n610), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n933), .A2(new_n722), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n220), .ZN(G1346gat));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n221), .B1(new_n933), .B2(new_n651), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n892), .A2(G162gat), .A3(new_n652), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n651), .B(new_n894), .C1(new_n920), .C2(new_n925), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G162gat), .ZN(new_n960));
  INV_X1    g759(.A(new_n957), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(KEYINPUT125), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n720), .A2(new_n434), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n865), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n266), .A3(new_n568), .ZN(new_n966));
  INV_X1    g765(.A(new_n965), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n723), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n266), .B2(new_n968), .ZN(G1348gat));
  NOR2_X1   g768(.A1(new_n965), .A2(new_n683), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(new_n267), .ZN(G1349gat));
  OAI21_X1  g770(.A(G183gat), .B1(new_n965), .B2(new_n880), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n610), .A2(new_n275), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT60), .ZN(G1350gat));
  OAI22_X1  g774(.A1(new_n965), .A2(new_n652), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(G1351gat));
  INV_X1    g777(.A(new_n889), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n720), .A2(new_n432), .A3(new_n434), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n723), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n948), .A2(new_n980), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n569), .A2(G197gat), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1352gat));
  OAI21_X1  g785(.A(G204gat), .B1(new_n983), .B2(new_n683), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n683), .A2(G204gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n979), .A2(new_n980), .A3(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n987), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1353gat));
  NAND3_X1  g795(.A1(new_n948), .A2(new_n610), .A3(new_n980), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G211gat), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT63), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(KEYINPUT127), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n728), .A2(G211gat), .ZN(new_n1005));
  AOI22_X1  g804(.A1(new_n1003), .A2(new_n1004), .B1(new_n981), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1002), .A2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(G218gat), .B1(new_n983), .B2(new_n652), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n981), .A2(new_n210), .A3(new_n651), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1355gat));
endmodule


