//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n207), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n210), .B(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n219), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  INV_X1    g0050(.A(new_n214), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n251), .A2(new_n252), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n258), .B1(G226), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n273), .A2(G223), .B1(new_n265), .B2(G77), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n262), .B1(new_n275), .B2(new_n259), .ZN(new_n276));
  INV_X1    g0076(.A(G190), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT69), .B(G200), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n254), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  XOR2_X1   g0083(.A(new_n283), .B(KEYINPUT66), .Z(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n214), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n287), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n284), .A2(new_n290), .B1(new_n202), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n214), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n203), .A2(KEYINPUT65), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n215), .A2(G33), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n294), .B1(new_n295), .B2(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT65), .B1(new_n203), .B2(G20), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n281), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n276), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n303), .B1(new_n310), .B2(G169), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n258), .B1(G244), .B2(new_n261), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n266), .A2(G232), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n273), .A2(G238), .B1(new_n265), .B2(G107), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(new_n259), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n277), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n280), .B2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n299), .A2(new_n297), .B1(new_n215), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n298), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n293), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT67), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n254), .B2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n290), .A2(new_n331), .B1(new_n324), .B2(new_n291), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(KEYINPUT68), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(KEYINPUT68), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n323), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n320), .A2(G179), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n320), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n335), .B2(new_n334), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n315), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n271), .A2(new_n272), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n226), .A2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(G226), .C2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n259), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n257), .B1(new_n260), .B2(new_n220), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n339), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT70), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n351), .A2(new_n352), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n353), .A2(new_n354), .B1(new_n360), .B2(new_n312), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n291), .A2(new_n219), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n290), .A2(G68), .A3(new_n282), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n297), .A2(new_n202), .B1(new_n215), .B2(G68), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n298), .A2(new_n324), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n293), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n365), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n369), .A2(new_n370), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n360), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G190), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n373), .C1(new_n378), .C2(new_n376), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n343), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n299), .B1(new_n254), .B2(G20), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n290), .A2(new_n382), .B1(new_n291), .B2(new_n299), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT71), .B1(new_n263), .B2(new_n264), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n271), .A2(new_n385), .A3(new_n272), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(new_n215), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n272), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n219), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n393), .B2(new_n201), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n296), .A2(G159), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT72), .B(G20), .C1(new_n393), .C2(new_n201), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n293), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n271), .A2(new_n215), .A3(new_n272), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n388), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT73), .A3(new_n390), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n265), .A2(new_n404), .A3(KEYINPUT7), .A4(new_n215), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(G68), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT16), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n383), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n257), .B1(new_n260), .B2(new_n226), .ZN(new_n410));
  INV_X1    g0210(.A(G226), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G1698), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n412), .B1(G223), .B2(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n259), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G179), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n339), .B2(new_n416), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n381), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n409), .A2(new_n381), .A3(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(new_n407), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n390), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n387), .B2(new_n388), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n407), .B(KEYINPUT16), .C1(new_n428), .C2(new_n219), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n293), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n413), .A2(new_n414), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n261), .A2(G232), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(new_n277), .A3(new_n257), .A4(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n378), .B1(new_n410), .B2(new_n415), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n430), .A2(KEYINPUT74), .A3(new_n383), .A4(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n383), .B(new_n437), .C1(new_n400), .C2(new_n408), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n423), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n423), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n422), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n380), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n289), .B1(new_n254), .B2(G33), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G107), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT25), .B1(new_n291), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n452), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n451), .A2(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT84), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n344), .A2(new_n215), .A3(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n344), .A2(new_n215), .A3(G87), .A4(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n215), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n452), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT24), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n464), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n458), .B1(new_n475), .B2(new_n293), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n464), .A2(new_n473), .A3(new_n470), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n464), .B2(new_n470), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n458), .B(new_n293), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n457), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n482));
  OAI211_X1 g0282(.A(G250), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G294), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n432), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  INV_X1    g0287(.A(G41), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT5), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(KEYINPUT79), .B2(G41), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n253), .A2(new_n489), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n493), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G264), .A3(new_n259), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n486), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n497), .A2(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(KEYINPUT85), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(G169), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n486), .A2(G179), .A3(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n494), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n481), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n293), .B1(new_n477), .B2(new_n478), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n456), .B1(new_n509), .B2(new_n479), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n378), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n498), .A2(new_n499), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(G190), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n215), .C1(G33), .C2(new_n227), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n293), .C1(new_n215), .C2(G116), .ZN(new_n518));
  XOR2_X1   g0318(.A(new_n518), .B(KEYINPUT20), .Z(new_n519));
  NOR2_X1   g0319(.A1(new_n287), .A2(G116), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n450), .B2(G116), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n271), .A2(G303), .A3(new_n272), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n524), .A2(new_n525), .A3(new_n529), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n432), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n495), .A2(G270), .A3(new_n259), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n494), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT81), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n494), .A2(new_n532), .A3(KEYINPUT81), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n523), .A2(new_n312), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n522), .A2(G169), .A3(new_n537), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n495), .A2(new_n259), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n494), .B1(new_n543), .B2(new_n228), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT4), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n516), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n273), .B2(G250), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n544), .B1(new_n553), .B2(new_n432), .ZN(new_n554));
  OR3_X1    g0354(.A1(new_n554), .A2(KEYINPUT80), .A3(new_n378), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT80), .B1(new_n554), .B2(new_n378), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n291), .A2(new_n227), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT77), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G97), .B2(new_n450), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n403), .A2(G107), .A3(new_n405), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n227), .A2(G107), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n452), .A2(G97), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n562), .B2(new_n563), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n566), .A2(new_n215), .B1(new_n324), .B2(new_n297), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n293), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n552), .A2(new_n550), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n549), .B1(new_n545), .B2(new_n546), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n432), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n544), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n277), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n554), .A2(new_n312), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n560), .A2(new_n568), .B1(new_n339), .B2(new_n574), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n557), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n522), .B1(G200), .B2(new_n537), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n277), .B2(new_n537), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n582));
  OAI211_X1 g0382(.A(G238), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n465), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n432), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n491), .A2(new_n222), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n253), .A2(new_n491), .B1(new_n586), .B2(new_n259), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n279), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n344), .A2(new_n215), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n215), .B1(new_n347), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n221), .A2(new_n227), .A3(new_n452), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n298), .B2(new_n227), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n293), .B1(new_n291), .B2(new_n326), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n451), .B2(new_n221), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n585), .A2(new_n587), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n277), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n589), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n597), .ZN(new_n602));
  INV_X1    g0402(.A(new_n326), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n450), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n339), .B1(new_n585), .B2(new_n587), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n312), .B2(new_n599), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n542), .A2(new_n579), .A3(new_n581), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n449), .A2(new_n515), .A3(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n379), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n361), .B1(new_n356), .B2(new_n358), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n341), .B1(new_n613), .B2(new_n373), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n438), .A2(new_n441), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n444), .B1(new_n615), .B2(KEYINPUT17), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n422), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n309), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n314), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT87), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n607), .B(new_n620), .C1(new_n312), .C2(new_n599), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n599), .A2(new_n312), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT87), .B1(new_n622), .B2(new_n606), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n604), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n601), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n578), .A2(new_n577), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n609), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n542), .ZN(new_n632));
  INV_X1    g0432(.A(new_n503), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n510), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n579), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n514), .A2(new_n625), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n629), .B(new_n631), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n619), .B1(new_n448), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT88), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n286), .A2(new_n215), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G213), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n632), .A2(new_n522), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n645), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n542), .B(new_n581), .C1(new_n523), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n515), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n510), .B2(new_n647), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n507), .B2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(new_n647), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n515), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n634), .B2(new_n647), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n208), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n593), .A2(G116), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G1), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n212), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT29), .B1(new_n637), .B2(new_n647), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n514), .A2(new_n625), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n507), .A2(new_n542), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n557), .A2(new_n576), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT92), .B1(new_n671), .B2(new_n627), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT92), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n579), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n669), .A2(new_n670), .A3(new_n672), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n624), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n628), .B1(new_n625), .B2(new_n627), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n645), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n668), .B1(KEYINPUT29), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n531), .A2(new_n535), .A3(new_n536), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n497), .A2(new_n312), .A3(new_n599), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n554), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n486), .A2(G179), .A3(new_n496), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n599), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n494), .A2(new_n532), .A3(KEYINPUT81), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT81), .B1(new_n494), .B2(new_n532), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n686), .A2(new_n554), .A3(new_n531), .A4(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT30), .B1(new_n690), .B2(KEYINPUT89), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n682), .A2(new_n692), .A3(new_n554), .A4(new_n686), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n684), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT91), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n501), .A2(new_n588), .A3(new_n572), .A4(new_n573), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT89), .B1(new_n698), .B2(new_n537), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n695), .A3(new_n693), .ZN(new_n700));
  INV_X1    g0500(.A(new_n684), .ZN(new_n701));
  AND4_X1   g0501(.A1(KEYINPUT91), .A2(new_n700), .A3(new_n696), .A4(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n645), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND4_X1   g0505(.A1(new_n542), .A2(new_n579), .A3(new_n581), .A4(new_n609), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n653), .A3(new_n647), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n647), .A2(new_n704), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n696), .B1(new_n694), .B2(KEYINPUT90), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n681), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n667), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n285), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n254), .B1(new_n716), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n662), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n652), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n650), .A2(new_n651), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n215), .A2(G179), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n279), .A2(new_n724), .A3(new_n277), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G87), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n215), .A2(new_n312), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n277), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT94), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n726), .B1(new_n734), .B2(new_n225), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G190), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n727), .A2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n277), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n344), .B1(new_n324), .B2(new_n737), .C1(new_n740), .C2(new_n202), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(G190), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G68), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n723), .A2(new_n736), .ZN(new_n744));
  INV_X1    g0544(.A(G159), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n744), .A2(KEYINPUT32), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT32), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n728), .A2(new_n312), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G97), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n743), .A2(new_n746), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n279), .A2(new_n724), .A3(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n452), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n735), .A2(new_n741), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n757));
  INV_X1    g0557(.A(new_n742), .ZN(new_n758));
  OR2_X1    g0558(.A1(KEYINPUT33), .A2(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(KEYINPUT33), .A2(G317), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(G294), .B2(new_n749), .ZN(new_n762));
  INV_X1    g0562(.A(G329), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n265), .B1(new_n744), .B2(new_n763), .C1(new_n764), .C2(new_n737), .ZN(new_n765));
  INV_X1    g0565(.A(new_n734), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(G322), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n739), .A2(G326), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G283), .A2(new_n752), .B1(new_n725), .B2(G303), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n762), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n757), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n214), .B1(G20), .B2(new_n339), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n661), .A2(new_n265), .ZN(new_n774));
  INV_X1    g0574(.A(G116), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G355), .A2(new_n774), .B1(new_n775), .B2(new_n661), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n384), .A2(new_n386), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n661), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n212), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n248), .A2(new_n490), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT93), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n781), .B2(new_n782), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n772), .A2(new_n773), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n784), .B(KEYINPUT96), .Z(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n649), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n722), .B1(new_n719), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT97), .ZN(G396));
  AND2_X1   g0592(.A1(new_n637), .A2(new_n647), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n335), .A2(new_n334), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(KEYINPUT102), .A3(new_n340), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT102), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n341), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n336), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n794), .A2(new_n645), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n336), .A2(new_n795), .A3(new_n801), .A4(new_n797), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n342), .A2(new_n645), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n713), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n719), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n773), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n719), .B1(G77), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n737), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n739), .A2(G137), .B1(new_n812), .B2(G159), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n295), .B2(new_n758), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G143), .B2(new_n766), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT100), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n752), .A2(G68), .ZN(new_n818));
  INV_X1    g0618(.A(new_n725), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n202), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n777), .B1(new_n822), .B2(new_n744), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n749), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n817), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n758), .A2(new_n827), .B1(new_n737), .B2(new_n775), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(KEYINPUT98), .B1(G303), .B2(new_n739), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(KEYINPUT98), .B2(new_n828), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT99), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n766), .A2(G294), .B1(G107), .B2(new_n725), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n752), .A2(G87), .ZN(new_n833));
  INV_X1    g0633(.A(new_n744), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n344), .B1(new_n834), .B2(G311), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n832), .A2(new_n750), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n825), .A2(new_n826), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n811), .B1(new_n837), .B2(new_n773), .ZN(new_n838));
  INV_X1    g0638(.A(new_n809), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n804), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n808), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(G116), .B(new_n216), .C1(new_n566), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n843), .B2(new_n566), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n213), .A2(G77), .A3(new_n392), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n254), .B(G13), .C1(new_n847), .C2(new_n244), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n610), .A2(new_n515), .A3(new_n645), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n708), .B1(new_n697), .B2(new_n702), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT108), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT91), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n700), .A2(new_n701), .ZN(new_n855));
  INV_X1    g0655(.A(new_n696), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n694), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(KEYINPUT108), .A3(new_n708), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n850), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n863), .A3(new_n645), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n864), .A3(new_n704), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n438), .A2(new_n441), .ZN(new_n867));
  INV_X1    g0667(.A(new_n391), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT16), .B1(new_n868), .B2(new_n407), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n383), .B1(new_n869), .B2(new_n400), .ZN(new_n870));
  INV_X1    g0670(.A(new_n643), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n418), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n409), .A2(new_n418), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n409), .A2(new_n871), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n873), .A2(KEYINPUT37), .B1(new_n867), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n871), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n409), .A2(new_n381), .A3(new_n418), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n419), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n880), .B(new_n881), .C1(new_n616), .C2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n883), .B(new_n443), .C1(new_n867), .C2(new_n423), .ZN(new_n885));
  INV_X1    g0685(.A(new_n881), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT104), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT38), .B(new_n879), .C1(new_n884), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n877), .B2(new_n867), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n445), .A2(new_n875), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n874), .A2(new_n875), .A3(new_n439), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n804), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n374), .A2(new_n645), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n379), .B(new_n896), .C1(new_n613), .C2(new_n373), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n374), .B(new_n645), .C1(new_n363), .C2(new_n612), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND4_X1   g0699(.A1(KEYINPUT40), .A2(new_n866), .A3(new_n894), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n804), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n865), .B2(new_n861), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n880), .B1(new_n445), .B2(new_n881), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n885), .A2(KEYINPUT104), .A3(new_n886), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n906), .B2(new_n879), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n908), .B(new_n878), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT105), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n879), .B1(new_n884), .B2(new_n887), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n908), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n913), .B2(new_n888), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n903), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n917), .A2(new_n448), .A3(new_n866), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n448), .B2(new_n866), .ZN(new_n919));
  OR3_X1    g0719(.A1(new_n918), .A2(new_n919), .A3(new_n651), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n910), .A2(new_n914), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n645), .B1(new_n795), .B2(new_n797), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n793), .B2(new_n799), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n901), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n921), .A2(new_n927), .B1(new_n883), .B2(new_n871), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n375), .A2(new_n645), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n913), .B2(new_n888), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n888), .A2(new_n931), .A3(new_n893), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT106), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT39), .B1(new_n907), .B2(new_n909), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n888), .A2(new_n893), .A3(new_n931), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n930), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n619), .B1(new_n681), .B2(new_n448), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n920), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n254), .B2(new_n716), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n920), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n849), .B1(new_n944), .B2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n569), .A2(new_n645), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n672), .A2(new_n674), .A3(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(new_n507), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n645), .B1(new_n949), .B2(new_n626), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n627), .A2(new_n645), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n658), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n950), .B1(KEYINPUT42), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n598), .A2(new_n645), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n625), .B(new_n624), .S(new_n956), .Z(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT109), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n954), .A2(new_n955), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n652), .A2(new_n655), .A3(new_n952), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n662), .B(new_n965), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n659), .A2(new_n952), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT111), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n659), .A2(new_n952), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT44), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n656), .ZN(new_n976));
  INV_X1    g0776(.A(new_n658), .ZN(new_n977));
  INV_X1    g0777(.A(new_n657), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n655), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n652), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n714), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n976), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n967), .B1(new_n983), .B2(new_n714), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n964), .B1(new_n984), .B2(new_n718), .ZN(new_n985));
  INV_X1    g0785(.A(new_n778), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n785), .B1(new_n208), .B2(new_n326), .C1(new_n986), .C2(new_n239), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n719), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n766), .A2(G150), .B1(G58), .B2(new_n725), .ZN(new_n989));
  INV_X1    g0789(.A(new_n749), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n758), .A2(new_n745), .B1(new_n990), .B2(new_n219), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G143), .B2(new_n739), .ZN(new_n992));
  INV_X1    g0792(.A(G137), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n344), .B1(new_n744), .B2(new_n993), .C1(new_n202), .C2(new_n737), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G77), .B2(new_n752), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G303), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n734), .A2(new_n997), .B1(new_n764), .B2(new_n740), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT112), .Z(new_n999));
  INV_X1    g0799(.A(G294), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n758), .A2(new_n1000), .B1(new_n990), .B2(new_n452), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT113), .B(G317), .Z(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n744), .B1(new_n737), .B2(new_n827), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1001), .A2(new_n777), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n752), .A2(G97), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT46), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n819), .B2(new_n775), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n725), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n996), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n988), .B1(new_n1011), .B2(new_n773), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n959), .B2(new_n789), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n985), .A2(new_n1013), .ZN(G387));
  OR2_X1    g0814(.A1(new_n655), .A2(new_n789), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n774), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1016), .A2(new_n664), .B1(G107), .B2(new_n208), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n986), .B1(new_n236), .B2(G45), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n664), .B(new_n490), .C1(new_n219), .C2(new_n324), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT114), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(KEYINPUT114), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT50), .B1(new_n299), .B2(G50), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n299), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1017), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n719), .B1(new_n1025), .B2(new_n786), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n734), .A2(new_n202), .B1(new_n324), .B2(new_n819), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n812), .A2(G68), .B1(new_n834), .B2(G150), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1028), .A2(new_n1005), .A3(new_n777), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n990), .A2(new_n326), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n299), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n742), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1030), .B(new_n1033), .C1(new_n745), .C2(new_n740), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n739), .A2(G322), .B1(new_n812), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n764), .B2(new_n758), .C1(new_n734), .C2(new_n1002), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n819), .A2(new_n1000), .B1(new_n827), .B2(new_n990), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n777), .B1(G326), .B2(new_n834), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n775), .B2(new_n753), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT115), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1026), .B1(new_n1047), .B2(new_n773), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n980), .A2(new_n718), .B1(new_n1015), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n981), .A2(new_n662), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n980), .A2(new_n714), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n976), .A2(new_n718), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n948), .A2(new_n784), .A3(new_n951), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n766), .A2(G311), .B1(G317), .B2(new_n739), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  AOI22_X1  g0857(.A1(G116), .A2(new_n749), .B1(new_n812), .B2(G294), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n997), .B2(new_n758), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT117), .Z(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n265), .B1(new_n744), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1062), .B(new_n754), .C1(G283), .C2(new_n725), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n734), .A2(new_n745), .B1(new_n295), .B2(new_n740), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n990), .A2(new_n324), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n834), .A2(G143), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n777), .C1(new_n299), .C2(new_n737), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G50), .C2(new_n742), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n725), .A2(G68), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n833), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n773), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n785), .B1(new_n227), .B2(new_n208), .C1(new_n986), .C2(new_n243), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1055), .A2(new_n719), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n983), .A2(new_n662), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n976), .A2(new_n982), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1053), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(G390));
  AOI21_X1  g0879(.A(new_n651), .B1(new_n861), .B2(new_n865), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n448), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n941), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT119), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n651), .B(new_n895), .C1(new_n861), .C2(new_n865), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n901), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n804), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n901), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(KEYINPUT119), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT118), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n645), .B(new_n798), .C1(new_n675), .C2(new_n679), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n922), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n680), .A2(new_n799), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n922), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(KEYINPUT118), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n712), .A2(G330), .A3(new_n804), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1091), .A2(new_n1094), .B1(new_n1095), .B2(new_n901), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1085), .A2(new_n1088), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1080), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n902), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1095), .A2(new_n901), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n926), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1082), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n930), .B1(new_n925), .B2(new_n1087), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n934), .A2(new_n938), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1091), .A2(new_n1094), .A3(new_n901), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n930), .A3(new_n894), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1095), .A2(new_n901), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1099), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1103), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1099), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n1102), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n662), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n934), .A2(new_n938), .A3(new_n809), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n719), .B1(new_n1032), .B2(new_n810), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n740), .A2(new_n1121), .B1(new_n990), .B2(new_n745), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G137), .B2(new_n742), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n344), .B1(new_n744), .B2(new_n1124), .C1(new_n737), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n766), .B2(G132), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1123), .B(new_n1127), .C1(new_n202), .C2(new_n753), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n725), .A2(G150), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1067), .B1(G107), .B2(new_n742), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n827), .B2(new_n740), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n766), .A2(G116), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n265), .B1(new_n737), .B2(new_n227), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G294), .B2(new_n834), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n726), .A3(new_n818), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1128), .A2(new_n1130), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1120), .B1(new_n1137), .B2(new_n773), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1118), .A2(new_n718), .B1(new_n1119), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1117), .A2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT122), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n928), .A2(new_n939), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n303), .A2(new_n871), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n315), .B(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n917), .B2(G330), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n894), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n866), .A2(new_n899), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT105), .B1(new_n907), .B2(new_n909), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n913), .A2(new_n911), .A3(new_n888), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n1148), .C1(new_n1152), .C2(KEYINPUT40), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1146), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1142), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n915), .A2(new_n916), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(G330), .A3(new_n1148), .A4(new_n1146), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n940), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1082), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1156), .A2(new_n1160), .B1(new_n1116), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1141), .B1(new_n1162), .B2(KEYINPUT57), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n663), .B1(new_n1162), .B2(KEYINPUT57), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n940), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n940), .B1(new_n1159), .B2(new_n1157), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1082), .B1(new_n1118), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT122), .B(new_n1165), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1163), .A2(new_n1164), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1168), .A2(new_n717), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1154), .A2(new_n809), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n719), .B1(G50), .B2(new_n810), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n758), .A2(new_n822), .B1(new_n740), .B2(new_n1124), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n990), .A2(new_n295), .B1(new_n737), .B2(new_n993), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1121), .B2(new_n734), .C1(new_n819), .C2(new_n1125), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n752), .A2(G159), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n834), .C2(G124), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n384), .A2(new_n386), .A3(new_n488), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n753), .A2(new_n225), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G107), .C2(new_n766), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n812), .A2(new_n603), .B1(new_n834), .B2(G283), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n227), .B2(new_n758), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G77), .B2(new_n725), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n739), .A2(G116), .B1(new_n749), .B2(G68), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT120), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1188), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT58), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1186), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1185), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1175), .B1(new_n1197), .B2(new_n773), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1173), .B1(new_n1174), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1172), .A2(new_n1199), .ZN(G375));
  NAND3_X1  g1000(.A1(new_n1097), .A2(new_n1101), .A3(new_n1082), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1103), .A2(new_n966), .A3(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(new_n1203));
  NAND2_X1  g1003(.A1(new_n1169), .A2(new_n718), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n719), .B1(G68), .B2(new_n810), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n734), .A2(new_n993), .B1(new_n745), .B2(new_n819), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n777), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n737), .A2(new_n295), .B1(new_n744), .B2(new_n1121), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1187), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n739), .A2(G132), .B1(new_n749), .B2(G50), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n758), .C2(new_n1125), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1031), .B1(G116), .B2(new_n742), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1000), .B2(new_n740), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n265), .B1(new_n744), .B2(new_n997), .C1(new_n452), .C2(new_n737), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G77), .B2(new_n752), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n227), .B2(new_n819), .C1(new_n827), .C2(new_n734), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1211), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1205), .B1(new_n1217), .B2(new_n773), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n901), .B2(new_n839), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1204), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1203), .A2(new_n1221), .ZN(G381));
  OR2_X1    g1022(.A1(G393), .A2(G396), .ZN(new_n1223));
  OR4_X1    g1023(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G381), .ZN(new_n1225));
  XOR2_X1   g1025(.A(G378), .B(KEYINPUT124), .Z(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(new_n1199), .A3(new_n1172), .A4(new_n1226), .ZN(G407));
  NAND2_X1  g1027(.A1(new_n644), .A2(G213), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G407), .B(G213), .C1(G375), .C2(new_n1230), .ZN(G409));
  NAND3_X1  g1031(.A1(new_n1172), .A2(G378), .A3(new_n1199), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1172), .A2(new_n1199), .A3(KEYINPUT125), .A4(G378), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1162), .A2(new_n966), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1199), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1226), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1228), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1169), .A2(new_n1242), .A3(new_n1161), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(new_n663), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1201), .B1(new_n1102), .B2(new_n1242), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G384), .B1(new_n1246), .B2(new_n1221), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n841), .B(new_n1220), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1229), .A2(G2897), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(G2897), .A3(new_n1229), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1254), .B2(new_n1250), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1241), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1240), .A2(new_n1228), .A3(new_n1249), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  XOR2_X1   g1059(.A(G393), .B(G396), .Z(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(G387), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1262), .A2(G390), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(G390), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G387), .B(G390), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1260), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1229), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1256), .A2(new_n1259), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(new_n1250), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1257), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1270), .A2(KEYINPUT62), .A3(new_n1249), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1268), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1265), .A2(new_n1267), .A3(KEYINPUT127), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1272), .B1(new_n1280), .B2(new_n1284), .ZN(G405));
  NAND2_X1  g1085(.A1(new_n1226), .A2(G375), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1236), .A2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1287), .A2(new_n1249), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1249), .ZN(new_n1289));
  OR3_X1    g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1268), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1268), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


