

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762;

  NOR2_X1 U381 ( .A1(n737), .A2(n742), .ZN(n738) );
  NOR2_X1 U382 ( .A1(n715), .A2(n710), .ZN(n645) );
  AND2_X1 U383 ( .A1(n745), .A2(KEYINPUT2), .ZN(n359) );
  OR2_X1 U384 ( .A1(n734), .A2(G902), .ZN(n400) );
  AND2_X1 U385 ( .A1(n370), .A2(n368), .ZN(n388) );
  INV_X1 U386 ( .A(n718), .ZN(n715) );
  INV_X2 U387 ( .A(n635), .ZN(n408) );
  NAND2_X2 U388 ( .A1(n568), .A2(n476), .ZN(n477) );
  NAND2_X2 U389 ( .A1(n389), .A2(n396), .ZN(n586) );
  AND2_X2 U390 ( .A1(n359), .A2(n688), .ZN(n635) );
  AND2_X2 U391 ( .A1(n392), .A2(n360), .ZN(n389) );
  AND2_X4 U392 ( .A1(n407), .A2(n408), .ZN(n733) );
  NOR2_X2 U393 ( .A1(n643), .A2(n509), .ZN(n510) );
  XNOR2_X2 U394 ( .A(n586), .B(KEYINPUT19), .ZN(n568) );
  XNOR2_X2 U395 ( .A(n514), .B(n513), .ZN(n516) );
  OR2_X2 U396 ( .A1(n699), .A2(n393), .ZN(n392) );
  INV_X1 U397 ( .A(n535), .ZN(n508) );
  AND2_X1 U398 ( .A1(n376), .A2(n506), .ZN(n507) );
  NOR2_X1 U399 ( .A1(n589), .A2(n588), .ZN(n724) );
  NOR2_X1 U400 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U401 ( .A(n380), .B(n379), .ZN(n639) );
  AND2_X1 U402 ( .A1(n392), .A2(n395), .ZN(n390) );
  XNOR2_X1 U403 ( .A(n501), .B(n743), .ZN(n734) );
  XNOR2_X1 U404 ( .A(n488), .B(n401), .ZN(n457) );
  XNOR2_X1 U405 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U406 ( .A(G137), .B(G146), .ZN(n441) );
  XNOR2_X1 U407 ( .A(KEYINPUT77), .B(G469), .ZN(n435) );
  INV_X1 U408 ( .A(G953), .ZN(n747) );
  OR2_X1 U409 ( .A1(n516), .A2(n649), .ZN(n529) );
  XNOR2_X1 U410 ( .A(n455), .B(n454), .ZN(n693) );
  NOR2_X2 U411 ( .A1(n632), .A2(n742), .ZN(n633) );
  XNOR2_X1 U412 ( .A(n457), .B(n430), .ZN(n438) );
  NOR2_X2 U413 ( .A1(n625), .A2(n624), .ZN(n745) );
  BUF_X1 U414 ( .A(n628), .Z(n688) );
  INV_X1 U415 ( .A(n438), .ZN(n383) );
  INV_X1 U416 ( .A(KEYINPUT10), .ZN(n413) );
  XOR2_X1 U417 ( .A(G137), .B(KEYINPUT74), .Z(n431) );
  XNOR2_X1 U418 ( .A(n429), .B(KEYINPUT25), .ZN(n367) );
  XOR2_X1 U419 ( .A(KEYINPUT83), .B(KEYINPUT5), .Z(n442) );
  XNOR2_X1 U420 ( .A(G131), .B(KEYINPUT84), .ZN(n444) );
  INV_X1 U421 ( .A(G237), .ZN(n465) );
  INV_X1 U422 ( .A(KEYINPUT8), .ZN(n415) );
  NAND2_X1 U423 ( .A1(n747), .A2(G234), .ZN(n416) );
  XNOR2_X1 U424 ( .A(KEYINPUT75), .B(G134), .ZN(n430) );
  XNOR2_X1 U425 ( .A(G134), .B(G122), .ZN(n484) );
  XOR2_X1 U426 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n482) );
  XNOR2_X1 U427 ( .A(n438), .B(n431), .ZN(n744) );
  XNOR2_X1 U428 ( .A(n411), .B(n374), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n375), .B(G104), .ZN(n374) );
  AND2_X1 U430 ( .A1(G227), .A2(n364), .ZN(n411) );
  INV_X1 U431 ( .A(G107), .ZN(n375) );
  XOR2_X1 U432 ( .A(KEYINPUT85), .B(G101), .Z(n433) );
  XNOR2_X1 U433 ( .A(G110), .B(G146), .ZN(n432) );
  NOR2_X1 U434 ( .A1(n589), .A2(n652), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n382), .B(KEYINPUT6), .ZN(n381) );
  INV_X1 U436 ( .A(KEYINPUT100), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n682), .B(n681), .ZN(n683) );
  XOR2_X1 U438 ( .A(n424), .B(n423), .Z(n630) );
  XNOR2_X1 U439 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U440 ( .A(n500), .B(n414), .ZN(n422) );
  XNOR2_X1 U441 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U442 ( .A1(n405), .A2(n361), .ZN(n407) );
  AND2_X1 U443 ( .A1(n631), .A2(G953), .ZN(n742) );
  INV_X1 U444 ( .A(KEYINPUT90), .ZN(n590) );
  XNOR2_X1 U445 ( .A(n365), .B(KEYINPUT103), .ZN(n541) );
  AND2_X1 U446 ( .A1(n759), .A2(n538), .ZN(n365) );
  NAND2_X1 U447 ( .A1(G237), .A2(G234), .ZN(n471) );
  INV_X1 U448 ( .A(G116), .ZN(n443) );
  XNOR2_X1 U449 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X1 U450 ( .A1(G953), .A2(G237), .ZN(n493) );
  INV_X1 U451 ( .A(KEYINPUT33), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n377), .A2(n649), .ZN(n380) );
  NAND2_X1 U453 ( .A1(n626), .A2(n467), .ZN(n395) );
  NAND2_X1 U454 ( .A1(n464), .A2(n394), .ZN(n393) );
  INV_X1 U455 ( .A(n467), .ZN(n394) );
  XNOR2_X1 U456 ( .A(KEYINPUT78), .B(KEYINPUT24), .ZN(n414) );
  XNOR2_X1 U457 ( .A(G128), .B(G119), .ZN(n417) );
  INV_X1 U458 ( .A(G122), .ZN(n453) );
  XNOR2_X1 U459 ( .A(G143), .B(G113), .ZN(n496) );
  INV_X1 U460 ( .A(KEYINPUT88), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n412), .B(G125), .ZN(n456) );
  XNOR2_X1 U462 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n459) );
  XNOR2_X1 U463 ( .A(n502), .B(n399), .ZN(n398) );
  INV_X1 U464 ( .A(G475), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n485), .B(KEYINPUT9), .ZN(n486) );
  XNOR2_X1 U466 ( .A(n744), .B(n371), .ZN(n729) );
  XNOR2_X1 U467 ( .A(n372), .B(n434), .ZN(n371) );
  XNOR2_X1 U468 ( .A(n373), .B(n499), .ZN(n372) );
  INV_X1 U469 ( .A(n556), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n369), .B(KEYINPUT104), .ZN(n368) );
  NOR2_X2 U471 ( .A1(n600), .A2(n569), .ZN(n716) );
  INV_X1 U472 ( .A(KEYINPUT68), .ZN(n363) );
  NOR2_X1 U473 ( .A1(n685), .A2(n742), .ZN(n687) );
  XOR2_X1 U474 ( .A(n734), .B(KEYINPUT59), .Z(n735) );
  NOR2_X1 U475 ( .A1(n702), .A2(n742), .ZN(n703) );
  XNOR2_X1 U476 ( .A(n558), .B(n381), .ZN(n583) );
  AND2_X1 U477 ( .A1(n395), .A2(n391), .ZN(n360) );
  XOR2_X1 U478 ( .A(n627), .B(KEYINPUT71), .Z(n361) );
  XNOR2_X1 U479 ( .A(n510), .B(KEYINPUT101), .ZN(n512) );
  NAND2_X1 U480 ( .A1(n508), .A2(n536), .ZN(n643) );
  XNOR2_X1 U481 ( .A(n494), .B(n410), .ZN(n498) );
  NOR2_X2 U482 ( .A1(n511), .A2(n512), .ZN(n514) );
  XNOR2_X2 U483 ( .A(n477), .B(KEYINPUT0), .ZN(n511) );
  XNOR2_X1 U484 ( .A(n387), .B(n363), .ZN(n362) );
  NOR2_X2 U485 ( .A1(n760), .A2(n678), .ZN(n517) );
  XNOR2_X1 U486 ( .A(n517), .B(KEYINPUT92), .ZN(n523) );
  NOR2_X2 U487 ( .A1(G902), .A2(n739), .ZN(n490) );
  XNOR2_X1 U488 ( .A(n545), .B(n544), .ZN(n628) );
  NOR2_X2 U489 ( .A1(n362), .A2(n515), .ZN(n678) );
  NOR2_X1 U490 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U491 ( .A1(n480), .A2(G217), .ZN(n481) );
  XNOR2_X2 U492 ( .A(n416), .B(n415), .ZN(n480) );
  BUF_X2 U493 ( .A(n747), .Z(n364) );
  XNOR2_X1 U494 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U495 ( .A(n456), .B(n413), .ZN(n500) );
  NAND2_X1 U496 ( .A1(n366), .A2(n565), .ZN(n567) );
  NAND2_X1 U497 ( .A1(n563), .A2(n564), .ZN(n366) );
  XNOR2_X2 U498 ( .A(n428), .B(n367), .ZN(n515) );
  NOR2_X1 U499 ( .A1(n516), .A2(n378), .ZN(n370) );
  XNOR2_X1 U500 ( .A(n758), .B(KEYINPUT72), .ZN(n376) );
  XNOR2_X2 U501 ( .A(n402), .B(n505), .ZN(n758) );
  NAND2_X1 U502 ( .A1(n650), .A2(n649), .ZN(n533) );
  XNOR2_X2 U503 ( .A(n566), .B(n437), .ZN(n649) );
  AND2_X2 U504 ( .A1(n650), .A2(n378), .ZN(n377) );
  INV_X1 U505 ( .A(n583), .ZN(n378) );
  XNOR2_X1 U506 ( .A(n384), .B(n383), .ZN(n682) );
  XNOR2_X1 U507 ( .A(n447), .B(n440), .ZN(n384) );
  XNOR2_X2 U508 ( .A(n386), .B(n385), .ZN(n452) );
  XNOR2_X2 U509 ( .A(G119), .B(KEYINPUT3), .ZN(n385) );
  XNOR2_X2 U510 ( .A(G113), .B(G101), .ZN(n386) );
  NOR2_X1 U511 ( .A1(n516), .A2(n397), .ZN(n387) );
  XNOR2_X2 U512 ( .A(n388), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U513 ( .A1(n396), .A2(n390), .ZN(n621) );
  INV_X1 U514 ( .A(n641), .ZN(n391) );
  NAND2_X1 U515 ( .A1(n699), .A2(n467), .ZN(n396) );
  NOR2_X2 U516 ( .A1(n639), .A2(n478), .ZN(n479) );
  OR2_X1 U517 ( .A1(n649), .A2(n559), .ZN(n397) );
  XNOR2_X2 U518 ( .A(n400), .B(n398), .ZN(n535) );
  XNOR2_X2 U519 ( .A(G143), .B(G128), .ZN(n488) );
  NAND2_X1 U520 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U521 ( .A(n479), .B(KEYINPUT34), .ZN(n404) );
  XNOR2_X1 U522 ( .A(n546), .B(n409), .ZN(n406) );
  NAND2_X1 U523 ( .A1(n406), .A2(n745), .ZN(n405) );
  NOR2_X2 U524 ( .A1(G902), .A2(n729), .ZN(n436) );
  AND2_X1 U525 ( .A1(n493), .A2(G214), .ZN(n410) );
  INV_X1 U526 ( .A(KEYINPUT46), .ZN(n605) );
  XNOR2_X1 U527 ( .A(n605), .B(KEYINPUT64), .ZN(n606) );
  INV_X1 U528 ( .A(KEYINPUT89), .ZN(n610) );
  XNOR2_X1 U529 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n613), .B(n612), .ZN(n625) );
  XNOR2_X1 U531 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U532 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U533 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U534 ( .A(n677), .B(n676), .ZN(G75) );
  XNOR2_X1 U535 ( .A(n431), .B(KEYINPUT23), .ZN(n424) );
  INV_X1 U536 ( .A(G146), .ZN(n412) );
  NAND2_X1 U537 ( .A1(G221), .A2(n480), .ZN(n420) );
  XOR2_X1 U538 ( .A(G140), .B(G110), .Z(n418) );
  XOR2_X1 U539 ( .A(n418), .B(n417), .Z(n419) );
  XNOR2_X1 U540 ( .A(G902), .B(KEYINPUT15), .ZN(n464) );
  NAND2_X1 U541 ( .A1(n464), .A2(G234), .ZN(n425) );
  XNOR2_X1 U542 ( .A(n425), .B(KEYINPUT20), .ZN(n427) );
  NAND2_X1 U543 ( .A1(G221), .A2(n427), .ZN(n426) );
  XNOR2_X1 U544 ( .A(KEYINPUT21), .B(n426), .ZN(n509) );
  INV_X1 U545 ( .A(n509), .ZN(n653) );
  NAND2_X1 U546 ( .A1(n427), .A2(G217), .ZN(n429) );
  NOR2_X1 U547 ( .A1(n630), .A2(G902), .ZN(n428) );
  AND2_X2 U548 ( .A1(n653), .A2(n515), .ZN(n650) );
  XNOR2_X1 U549 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U550 ( .A(G140), .B(G131), .Z(n499) );
  XNOR2_X2 U551 ( .A(n436), .B(n435), .ZN(n566) );
  XNOR2_X1 U552 ( .A(KEYINPUT70), .B(KEYINPUT1), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n493), .A2(G210), .ZN(n439) );
  XNOR2_X1 U554 ( .A(n452), .B(n439), .ZN(n440) );
  XNOR2_X1 U555 ( .A(n442), .B(n441), .ZN(n446) );
  INV_X1 U556 ( .A(G902), .ZN(n466) );
  NAND2_X1 U557 ( .A1(n682), .A2(n466), .ZN(n449) );
  INV_X1 U558 ( .A(G472), .ZN(n448) );
  XNOR2_X2 U559 ( .A(n449), .B(n448), .ZN(n558) );
  XNOR2_X1 U560 ( .A(KEYINPUT79), .B(KEYINPUT16), .ZN(n450) );
  XNOR2_X1 U561 ( .A(n450), .B(G110), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n453), .B(G104), .ZN(n495) );
  XNOR2_X2 U564 ( .A(G116), .B(G107), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n495), .B(n483), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n457), .B(n456), .ZN(n462) );
  NAND2_X1 U567 ( .A1(n747), .A2(G224), .ZN(n458) );
  XNOR2_X1 U568 ( .A(n458), .B(KEYINPUT93), .ZN(n460) );
  XNOR2_X1 U569 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U571 ( .A(n463), .B(n693), .ZN(n699) );
  INV_X1 U572 ( .A(n464), .ZN(n626) );
  NAND2_X1 U573 ( .A1(n466), .A2(n465), .ZN(n468) );
  NAND2_X1 U574 ( .A1(n468), .A2(G210), .ZN(n467) );
  NAND2_X1 U575 ( .A1(n468), .A2(G214), .ZN(n470) );
  INV_X1 U576 ( .A(KEYINPUT94), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n470), .B(n469), .ZN(n641) );
  XNOR2_X1 U578 ( .A(KEYINPUT14), .B(n471), .ZN(n472) );
  NAND2_X1 U579 ( .A1(G952), .A2(n472), .ZN(n667) );
  NOR2_X1 U580 ( .A1(G953), .A2(n667), .ZN(n550) );
  NAND2_X1 U581 ( .A1(n472), .A2(G902), .ZN(n548) );
  OR2_X1 U582 ( .A1(n364), .A2(G898), .ZN(n694) );
  NOR2_X1 U583 ( .A1(n548), .A2(n694), .ZN(n473) );
  OR2_X1 U584 ( .A1(n550), .A2(n473), .ZN(n475) );
  INV_X1 U585 ( .A(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U586 ( .A(n475), .B(n474), .ZN(n476) );
  BUF_X1 U587 ( .A(n511), .Z(n478) );
  INV_X1 U588 ( .A(n478), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n482), .B(n481), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n489), .B(n488), .ZN(n739) );
  XNOR2_X2 U592 ( .A(G478), .B(n490), .ZN(n536) );
  INV_X1 U593 ( .A(n536), .ZN(n503) );
  XNOR2_X1 U594 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n502) );
  XOR2_X1 U595 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n492) );
  XNOR2_X1 U596 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n743) );
  NAND2_X1 U600 ( .A1(n503), .A2(n535), .ZN(n504) );
  XOR2_X1 U601 ( .A(KEYINPUT105), .B(n504), .Z(n556) );
  INV_X1 U602 ( .A(KEYINPUT35), .ZN(n505) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n506) );
  NOR2_X1 U604 ( .A1(n507), .A2(KEYINPUT67), .ZN(n521) );
  XNOR2_X1 U605 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n513) );
  BUF_X1 U606 ( .A(n515), .Z(n652) );
  INV_X1 U607 ( .A(n649), .ZN(n589) );
  AND2_X1 U608 ( .A1(n758), .A2(KEYINPUT72), .ZN(n518) );
  NAND2_X1 U609 ( .A1(n523), .A2(n518), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n519), .A2(KEYINPUT44), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n521), .A2(n520), .ZN(n527) );
  NAND2_X1 U612 ( .A1(n758), .A2(KEYINPUT67), .ZN(n522) );
  NAND2_X1 U613 ( .A1(n522), .A2(KEYINPUT44), .ZN(n525) );
  INV_X1 U614 ( .A(n523), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U616 ( .A1(n527), .A2(n526), .ZN(n543) );
  NAND2_X1 U617 ( .A1(n583), .A2(n652), .ZN(n528) );
  XOR2_X1 U618 ( .A(KEYINPUT102), .B(n530), .Z(n759) );
  NAND2_X1 U619 ( .A1(n566), .A2(n650), .ZN(n547) );
  NOR2_X1 U620 ( .A1(n547), .A2(n559), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n532), .A2(n531), .ZN(n707) );
  OR2_X1 U622 ( .A1(n533), .A2(n558), .ZN(n658) );
  NOR2_X1 U623 ( .A1(n658), .A2(n478), .ZN(n534) );
  XNOR2_X1 U624 ( .A(n534), .B(KEYINPUT31), .ZN(n720) );
  NAND2_X1 U625 ( .A1(n707), .A2(n720), .ZN(n537) );
  NAND2_X1 U626 ( .A1(n536), .A2(n535), .ZN(n718) );
  NOR2_X1 U627 ( .A1(n536), .A2(n535), .ZN(n710) );
  XOR2_X1 U628 ( .A(KEYINPUT86), .B(n645), .Z(n572) );
  NAND2_X1 U629 ( .A1(n537), .A2(n572), .ZN(n538) );
  INV_X1 U630 ( .A(KEYINPUT67), .ZN(n539) );
  NOR2_X1 U631 ( .A1(n539), .A2(KEYINPUT44), .ZN(n540) );
  NOR2_X1 U632 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U634 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n544) );
  NAND2_X1 U635 ( .A1(n628), .A2(n626), .ZN(n546) );
  INV_X1 U636 ( .A(n547), .ZN(n555) );
  OR2_X1 U637 ( .A1(n364), .A2(n548), .ZN(n549) );
  NOR2_X1 U638 ( .A1(G900), .A2(n549), .ZN(n551) );
  NOR2_X1 U639 ( .A1(n551), .A2(n550), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n641), .A2(n558), .ZN(n552) );
  XOR2_X1 U641 ( .A(KEYINPUT30), .B(n552), .Z(n553) );
  NOR2_X1 U642 ( .A1(n580), .A2(n553), .ZN(n554) );
  NAND2_X1 U643 ( .A1(n555), .A2(n554), .ZN(n594) );
  OR2_X1 U644 ( .A1(n594), .A2(n621), .ZN(n557) );
  NOR2_X1 U645 ( .A1(n557), .A2(n556), .ZN(n714) );
  INV_X1 U646 ( .A(n558), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n559), .A2(n653), .ZN(n560) );
  OR2_X1 U648 ( .A1(n580), .A2(n560), .ZN(n561) );
  NOR2_X1 U649 ( .A1(n652), .A2(n561), .ZN(n562) );
  NAND2_X1 U650 ( .A1(KEYINPUT28), .A2(n562), .ZN(n565) );
  INV_X1 U651 ( .A(KEYINPUT28), .ZN(n564) );
  INV_X1 U652 ( .A(n562), .ZN(n563) );
  NAND2_X1 U653 ( .A1(n567), .A2(n566), .ZN(n600) );
  INV_X1 U654 ( .A(n568), .ZN(n569) );
  INV_X1 U655 ( .A(n645), .ZN(n570) );
  NAND2_X1 U656 ( .A1(n716), .A2(n570), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n571), .A2(KEYINPUT47), .ZN(n577) );
  XNOR2_X1 U658 ( .A(KEYINPUT47), .B(KEYINPUT73), .ZN(n573) );
  NAND2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U660 ( .A(KEYINPUT81), .B(n574), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n716), .A2(n575), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U663 ( .A1(n714), .A2(n578), .ZN(n579) );
  XNOR2_X1 U664 ( .A(KEYINPUT80), .B(n579), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n580), .A2(n652), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n581), .A2(n653), .ZN(n582) );
  NOR2_X1 U667 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n584), .B(KEYINPUT106), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n585), .A2(n715), .ZN(n615) );
  NOR2_X1 U670 ( .A1(n615), .A2(n586), .ZN(n587) );
  XOR2_X1 U671 ( .A(KEYINPUT36), .B(n587), .Z(n588) );
  XNOR2_X1 U672 ( .A(n724), .B(n590), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n609) );
  XOR2_X1 U674 ( .A(KEYINPUT82), .B(KEYINPUT38), .Z(n593) );
  XNOR2_X1 U675 ( .A(n621), .B(n593), .ZN(n640) );
  NOR2_X1 U676 ( .A1(n640), .A2(n594), .ZN(n596) );
  XOR2_X1 U677 ( .A(KEYINPUT91), .B(KEYINPUT39), .Z(n595) );
  XNOR2_X1 U678 ( .A(n596), .B(n595), .ZN(n614) );
  NOR2_X1 U679 ( .A1(n718), .A2(n614), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n597), .B(KEYINPUT40), .ZN(n762) );
  INV_X1 U681 ( .A(KEYINPUT111), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n641), .A2(n640), .ZN(n598) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT109), .ZN(n644) );
  NOR2_X1 U684 ( .A1(n644), .A2(n643), .ZN(n599) );
  XNOR2_X1 U685 ( .A(n599), .B(KEYINPUT41), .ZN(n668) );
  NOR2_X1 U686 ( .A1(n668), .A2(n600), .ZN(n602) );
  XNOR2_X1 U687 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n601) );
  XNOR2_X1 U688 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n604), .B(n603), .ZN(n757) );
  NOR2_X1 U690 ( .A1(n762), .A2(n757), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(n606), .ZN(n608) );
  XOR2_X1 U692 ( .A(KEYINPUT76), .B(KEYINPUT48), .Z(n611) );
  INV_X1 U693 ( .A(n710), .ZN(n721) );
  NOR2_X1 U694 ( .A1(n614), .A2(n721), .ZN(n726) );
  INV_X1 U695 ( .A(n726), .ZN(n623) );
  INV_X1 U696 ( .A(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n641), .A2(n649), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U699 ( .A(KEYINPUT43), .B(n618), .ZN(n620) );
  XOR2_X1 U700 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n619) );
  XNOR2_X1 U701 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n680) );
  NAND2_X1 U703 ( .A1(n623), .A2(n680), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n733), .A2(G217), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(n630), .ZN(n632) );
  INV_X1 U707 ( .A(G952), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT122), .ZN(G66) );
  NOR2_X1 U709 ( .A1(n688), .A2(KEYINPUT2), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n745), .A2(KEYINPUT2), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT87), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n673) );
  BUF_X1 U714 ( .A(n639), .Z(n669) );
  AND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n669), .A2(n648), .ZN(n664) );
  OR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(KEYINPUT50), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U723 ( .A(KEYINPUT49), .B(n654), .Z(n655) );
  NOR2_X1 U724 ( .A1(n559), .A2(n655), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n661) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n662), .A2(n668), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT52), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U736 ( .A(KEYINPUT120), .B(n674), .Z(n675) );
  NAND2_X1 U737 ( .A1(n364), .A2(n675), .ZN(n677) );
  XNOR2_X1 U738 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n676) );
  XOR2_X1 U739 ( .A(n678), .B(G110), .Z(G12) );
  XNOR2_X1 U740 ( .A(G140), .B(KEYINPUT118), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n680), .B(n679), .ZN(G42) );
  NAND2_X1 U742 ( .A1(n733), .A2(G472), .ZN(n684) );
  XOR2_X1 U743 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n681) );
  XNOR2_X1 U744 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U745 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n687), .B(n686), .ZN(G57) );
  NAND2_X1 U747 ( .A1(n688), .A2(n364), .ZN(n692) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n689) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n689), .ZN(n690) );
  NAND2_X1 U750 ( .A1(n690), .A2(G898), .ZN(n691) );
  NAND2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U752 ( .A(n694), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n693), .A2(n695), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n697), .B(n696), .ZN(G69) );
  NAND2_X1 U755 ( .A1(n733), .A2(G210), .ZN(n701) );
  XOR2_X1 U756 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n698) );
  XNOR2_X1 U757 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U760 ( .A1(n718), .A2(n707), .ZN(n704) );
  XOR2_X1 U761 ( .A(G104), .B(n704), .Z(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n706) );
  XNOR2_X1 U763 ( .A(G107), .B(KEYINPUT27), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n706), .B(n705), .ZN(n709) );
  NOR2_X1 U765 ( .A1(n721), .A2(n707), .ZN(n708) );
  XOR2_X1 U766 ( .A(n709), .B(n708), .Z(G9) );
  XOR2_X1 U767 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n712) );
  NAND2_X1 U768 ( .A1(n716), .A2(n710), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U770 ( .A(G128), .B(n713), .Z(G30) );
  XOR2_X1 U771 ( .A(G143), .B(n714), .Z(G45) );
  NAND2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n717), .B(G146), .ZN(G48) );
  NOR2_X1 U774 ( .A1(n718), .A2(n720), .ZN(n719) );
  XOR2_X1 U775 ( .A(G113), .B(n719), .Z(G15) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U777 ( .A(KEYINPUT116), .B(n722), .Z(n723) );
  XNOR2_X1 U778 ( .A(G116), .B(n723), .ZN(G18) );
  XNOR2_X1 U779 ( .A(G125), .B(n724), .ZN(n725) );
  XNOR2_X1 U780 ( .A(n725), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U781 ( .A(G134), .B(n726), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n727), .B(KEYINPUT117), .ZN(G36) );
  NAND2_X1 U783 ( .A1(n733), .A2(G469), .ZN(n731) );
  XOR2_X1 U784 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n742), .A2(n732), .ZN(G54) );
  NAND2_X1 U787 ( .A1(n733), .A2(G475), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U790 ( .A1(n733), .A2(G478), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(G63) );
  XOR2_X1 U793 ( .A(n744), .B(n743), .Z(n750) );
  XOR2_X1 U794 ( .A(n745), .B(n750), .Z(n746) );
  XNOR2_X1 U795 ( .A(n746), .B(KEYINPUT123), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n364), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT124), .ZN(n756) );
  XNOR2_X1 U798 ( .A(G227), .B(KEYINPUT125), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U800 ( .A1(G900), .A2(n752), .ZN(n753) );
  XNOR2_X1 U801 ( .A(KEYINPUT126), .B(n753), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U804 ( .A(n757), .B(G137), .Z(G39) );
  XNOR2_X1 U805 ( .A(n758), .B(G122), .ZN(G24) );
  XNOR2_X1 U806 ( .A(G101), .B(n759), .ZN(G3) );
  XNOR2_X1 U807 ( .A(G119), .B(KEYINPUT127), .ZN(n761) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(G21) );
  XOR2_X1 U809 ( .A(G131), .B(n762), .Z(G33) );
endmodule

