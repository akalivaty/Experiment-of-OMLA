//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT64), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n215), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT8), .A2(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT67), .B(G58), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(KEYINPUT8), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n250), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n249), .B1(new_n206), .B2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(G50), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(new_n259), .B2(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n276), .A2(G223), .B1(G77), .B2(new_n274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n274), .A2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n254), .C2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(G226), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n282), .A2(new_n283), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n283), .B1(new_n282), .B2(new_n290), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n270), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n282), .A2(new_n290), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n282), .A2(new_n283), .A3(new_n290), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G200), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT10), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n298), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(G190), .B1(new_n268), .B2(new_n269), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n300), .A4(new_n299), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT12), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n219), .B1(new_n308), .B2(KEYINPUT70), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n262), .ZN(new_n311));
  INV_X1    g0111(.A(new_n262), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n312), .A2(KEYINPUT70), .A3(new_n308), .A4(new_n219), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n311), .A2(new_n313), .B1(new_n260), .B2(G68), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n255), .A2(G77), .B1(G20), .B2(new_n219), .ZN(new_n315));
  INV_X1    g0115(.A(new_n257), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n202), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n317), .A2(new_n318), .A3(new_n249), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n317), .B2(new_n249), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(KEYINPUT71), .B(new_n314), .C1(new_n319), .C2(new_n320), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT3), .B(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G232), .A3(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G226), .A3(new_n275), .ZN(new_n329));
  INV_X1    g0129(.A(G97), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n328), .B(new_n329), .C1(new_n254), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n281), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n286), .B1(G238), .B2(new_n289), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n332), .B2(new_n333), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n326), .B(G169), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n337), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G179), .A3(new_n335), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n335), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n326), .B1(new_n342), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n325), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n336), .A2(new_n337), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G190), .B1(new_n323), .B2(new_n324), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT69), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n342), .B2(G200), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n347), .B(G200), .C1(new_n336), .C2(new_n337), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n327), .A2(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G107), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n353), .A2(new_n220), .B1(new_n354), .B2(new_n327), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n274), .A2(new_n231), .A3(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n281), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n286), .B1(G244), .B2(new_n289), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n294), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT8), .B(G58), .Z(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n207), .A2(G33), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n249), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n260), .A2(G77), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(G77), .C2(new_n262), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n359), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n359), .A2(G179), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n368), .B1(new_n370), .B2(G169), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n369), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n293), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n264), .B1(new_n303), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n307), .A2(new_n352), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  MUX2_X1   g0182(.A(new_n312), .B(new_n260), .S(new_n253), .Z(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n201), .B1(new_n252), .B2(G68), .ZN(new_n385));
  INV_X1    g0185(.A(G159), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n385), .A2(new_n207), .B1(new_n386), .B2(new_n316), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n272), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n389));
  OAI211_X1 g0189(.A(KEYINPUT7), .B(new_n207), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n274), .A2(KEYINPUT72), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n327), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n387), .B1(new_n396), .B2(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT73), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n395), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n271), .B2(new_n273), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT72), .B1(new_n400), .B2(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT67), .A2(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT67), .A2(G58), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G58), .B2(G68), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n407));
  AND4_X1   g0207(.A1(KEYINPUT73), .A2(new_n402), .A3(KEYINPUT16), .A4(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n219), .B1(new_n395), .B2(new_n390), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT74), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n249), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n384), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n289), .A2(G232), .ZN(new_n420));
  INV_X1    g0220(.A(new_n286), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n278), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n276), .A2(G226), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n281), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n376), .B2(new_n426), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(new_n419), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n397), .A2(KEYINPUT73), .A3(KEYINPUT16), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n327), .A2(new_n394), .A3(G20), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT7), .B1(new_n274), .B2(new_n207), .ZN(new_n436));
  OAI21_X1  g0236(.A(G68), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT74), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n407), .A3(new_n413), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n250), .B1(new_n439), .B2(new_n410), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n383), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n428), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT18), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n429), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n426), .A2(new_n294), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G200), .B2(new_n426), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n384), .B(new_n446), .C1(new_n409), .C2(new_n417), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(KEYINPUT17), .A3(new_n446), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n381), .A2(new_n382), .A3(new_n444), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n307), .A2(new_n352), .A3(new_n380), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n429), .A2(new_n449), .A3(new_n443), .A4(new_n450), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT75), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n207), .C1(G33), .C2(new_n330), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n249), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n249), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n262), .A2(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  AND4_X1   g0268(.A1(new_n215), .A2(new_n262), .A3(new_n248), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(G116), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n466), .B1(new_n465), .B2(new_n470), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n281), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G270), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n477), .A2(new_n288), .A3(G274), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n327), .A2(G257), .A3(new_n275), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n274), .A2(G303), .ZN(new_n484));
  INV_X1    g0284(.A(G264), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n484), .C1(new_n353), .C2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n486), .A2(KEYINPUT79), .A3(new_n281), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT79), .B1(new_n486), .B2(new_n281), .ZN(new_n488));
  OAI211_X1 g0288(.A(G190), .B(new_n482), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n488), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(KEYINPUT79), .A3(new_n281), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n481), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n474), .B(new_n489), .C1(new_n492), .C2(new_n371), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  OAI21_X1  g0294(.A(G169), .B1(new_n472), .B2(new_n473), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n492), .ZN(new_n496));
  OAI211_X1 g0296(.A(G179), .B(new_n482), .C1(new_n487), .C2(new_n488), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n473), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n471), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT21), .A4(G169), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n493), .A2(new_n496), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n502), .A3(G169), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n503), .A4(new_n493), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n271), .A2(new_n273), .A3(G238), .A4(new_n275), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n281), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n281), .A2(new_n284), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n476), .A2(new_n222), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n516), .A2(new_n476), .B1(new_n288), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G200), .ZN(new_n520));
  INV_X1    g0320(.A(new_n364), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n262), .ZN(new_n522));
  NAND3_X1  g0322(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n207), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G97), .A2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n221), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n271), .A2(new_n273), .A3(new_n207), .A4(G68), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n363), .B2(new_n330), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n250), .B1(new_n531), .B2(KEYINPUT77), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT77), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n527), .A2(new_n528), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n522), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n250), .A2(new_n262), .A3(new_n468), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n221), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n520), .A2(new_n535), .A3(KEYINPUT78), .A4(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n515), .A2(new_n518), .A3(G190), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n522), .B(new_n537), .C1(new_n532), .C2(new_n534), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT78), .B1(new_n542), .B2(new_n520), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n532), .A2(new_n534), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n469), .A2(new_n521), .ZN(new_n546));
  INV_X1    g0346(.A(new_n522), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n515), .A2(new_n518), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n378), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n519), .A2(new_n376), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n271), .A2(new_n273), .A3(new_n207), .A4(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n327), .A2(new_n557), .A3(new_n207), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT82), .B1(new_n207), .B2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT23), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT82), .B(new_n563), .C1(new_n207), .C2(G107), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n562), .A2(new_n564), .B1(G116), .B2(new_n255), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n559), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n249), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT83), .B(new_n249), .C1(new_n566), .C2(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n354), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT25), .B1(new_n312), .B2(new_n354), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(new_n575), .B1(new_n536), .B2(new_n354), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n327), .A2(G257), .A3(G1698), .ZN(new_n579));
  INV_X1    g0379(.A(G294), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n327), .A2(new_n275), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n579), .B1(new_n254), .B2(new_n580), .C1(new_n581), .C2(new_n222), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n281), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n478), .A2(G264), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n480), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n376), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n582), .A2(new_n281), .B1(G264), .B2(new_n478), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n378), .A3(new_n480), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n578), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT6), .ZN(new_n592));
  AND2_X1   g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n525), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n354), .A2(KEYINPUT6), .A3(G97), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G77), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n596), .A2(new_n207), .B1(new_n597), .B2(new_n316), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n354), .B1(new_n395), .B2(new_n390), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n249), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n262), .A2(G97), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n469), .B2(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(KEYINPUT5), .A2(G41), .ZN(new_n604));
  NOR2_X1   g0404(.A1(KEYINPUT5), .A2(G41), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n476), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G257), .A3(new_n288), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n480), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(new_n275), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n327), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n327), .A2(G250), .A3(G1698), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n457), .A4(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n608), .B1(new_n614), .B2(new_n281), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n378), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n603), .B(new_n616), .C1(G169), .C2(new_n615), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT76), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(KEYINPUT76), .B(new_n608), .C1(new_n614), .C2(new_n281), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n615), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n600), .B(new_n602), .C1(new_n622), .C2(new_n294), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n617), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n576), .B1(new_n570), .B2(new_n571), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n585), .A2(new_n371), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G190), .B2(new_n585), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n591), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n456), .A2(new_n510), .A3(new_n554), .A4(new_n630), .ZN(G372));
  NAND4_X1  g0431(.A1(new_n520), .A2(new_n535), .A3(new_n538), .A4(new_n540), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n552), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n626), .B2(new_n628), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n496), .A2(new_n501), .A3(new_n503), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n589), .B1(new_n572), .B2(new_n577), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n634), .B(new_n625), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(G107), .B1(new_n435), .B2(new_n436), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n594), .A2(new_n595), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n250), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n602), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n615), .B2(G169), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n615), .A2(new_n378), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n645), .B(new_n552), .C1(new_n541), .C2(new_n543), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT26), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n633), .A2(new_n617), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n553), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n637), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n456), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n307), .B(KEYINPUT84), .ZN(new_n653));
  INV_X1    g0453(.A(new_n344), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n374), .A2(new_n373), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n351), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n451), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n444), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n653), .A2(new_n658), .B1(new_n377), .B2(new_n379), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n500), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n507), .B2(new_n503), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n510), .B2(new_n667), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n591), .A2(new_n629), .ZN(new_n672));
  INV_X1    g0472(.A(new_n666), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n626), .A2(new_n673), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n672), .A2(new_n674), .B1(new_n591), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n635), .A2(new_n673), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n672), .A2(new_n677), .B1(new_n591), .B2(new_n666), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n526), .A2(G116), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT85), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n213), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n510), .A2(new_n630), .A3(new_n554), .A4(new_n673), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n587), .A2(new_n549), .A3(new_n615), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n497), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(KEYINPUT30), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n549), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n502), .A2(new_n585), .A3(new_n622), .A4(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n691), .B2(KEYINPUT30), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n666), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n698), .B(new_n666), .C1(new_n692), .C2(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n670), .B1(new_n689), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n651), .A2(new_n673), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n646), .A2(new_n649), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n624), .A2(KEYINPUT86), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT86), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n617), .B(new_n710), .C1(new_n621), .C2(new_n623), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n707), .B(new_n552), .C1(new_n708), .C2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n701), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n688), .B1(new_n715), .B2(G1), .ZN(G364));
  INV_X1    g0516(.A(G13), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G45), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT87), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT87), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n682), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n669), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n215), .B1(G20), .B2(new_n376), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n681), .A2(new_n327), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n214), .A2(new_n475), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(new_n246), .C2(new_n475), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n681), .A2(new_n274), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n459), .B2(new_n681), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n731), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n207), .A2(G190), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT88), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n371), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(KEYINPUT88), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G283), .A2(new_n743), .B1(new_n746), .B2(G329), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n294), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n378), .A2(new_n371), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n749), .A2(new_n738), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G326), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n378), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n738), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G322), .A2(new_n756), .B1(new_n758), .B2(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n748), .A2(new_n740), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n274), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n744), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G294), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n747), .A2(new_n753), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n327), .B1(new_n221), .B2(new_n760), .C1(new_n742), .C2(new_n354), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT89), .ZN(new_n768));
  INV_X1    g0568(.A(new_n750), .ZN(new_n769));
  INV_X1    g0569(.A(new_n751), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n202), .B1(new_n770), .B2(new_n219), .ZN(new_n771));
  INV_X1    g0571(.A(new_n252), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n772), .A2(new_n755), .B1(new_n757), .B2(new_n597), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OR3_X1    g0574(.A1(new_n745), .A2(KEYINPUT32), .A3(new_n386), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT32), .B1(new_n745), .B2(new_n386), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n764), .A2(G97), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n766), .B1(new_n768), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n737), .B1(new_n779), .B2(new_n729), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n724), .B1(new_n728), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n669), .B(new_n670), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n724), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT90), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NOR2_X1   g0585(.A1(new_n729), .A2(new_n725), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n724), .B1(new_n597), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n729), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n221), .A2(new_n742), .B1(new_n745), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n274), .B(new_n777), .C1(new_n769), .C2(new_n761), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n770), .A2(new_n792), .B1(new_n580), .B2(new_n755), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n760), .A2(new_n354), .B1(new_n757), .B2(new_n459), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n790), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G143), .A2(new_n756), .B1(new_n758), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G137), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n769), .C1(new_n798), .C2(new_n770), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n327), .B1(new_n760), .B2(new_n202), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n252), .B2(new_n764), .ZN(new_n804));
  INV_X1    g0604(.A(G132), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n219), .B2(new_n742), .C1(new_n805), .C2(new_n745), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n795), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n368), .A2(new_n666), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n369), .B2(new_n372), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n373), .B2(new_n374), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n655), .A2(new_n673), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n787), .B1(new_n788), .B2(new_n808), .C1(new_n814), .C2(new_n726), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n651), .A2(new_n814), .A3(new_n673), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT92), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n702), .A2(new_n813), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n701), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n724), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n815), .B1(new_n822), .B2(new_n823), .ZN(G384));
  NOR2_X1   g0624(.A1(new_n718), .A2(new_n206), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n325), .A2(new_n666), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n344), .A2(new_n351), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT93), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT93), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n351), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n341), .A2(new_n343), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n325), .B(new_n666), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n813), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n689), .A2(new_n700), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n664), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n249), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n432), .B2(new_n433), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n840), .B2(new_n383), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n454), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n428), .B1(new_n840), .B2(new_n383), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n844), .A3(new_n447), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n418), .A2(new_n428), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n664), .B(KEYINPUT94), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n418), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n849), .A3(new_n850), .A4(new_n447), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n843), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n843), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT95), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n843), .A2(new_n852), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT95), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n843), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n837), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT96), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n447), .B1(new_n441), .B2(new_n442), .ZN(new_n867));
  INV_X1    g0667(.A(new_n848), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n441), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n851), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n454), .A2(new_n869), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n857), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n843), .A2(new_n852), .A3(KEYINPUT96), .A4(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n866), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n835), .A2(KEYINPUT40), .A3(new_n836), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n863), .A2(new_n864), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT98), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n456), .A2(new_n836), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(G330), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n816), .A2(new_n812), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n831), .A2(new_n834), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n855), .B2(new_n861), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n444), .A2(new_n848), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n654), .A2(new_n673), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n866), .A2(new_n874), .A3(new_n891), .A4(new_n875), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n853), .B2(new_n854), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n456), .A2(new_n704), .A3(new_n714), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n659), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n825), .B1(new_n883), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n883), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n639), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n639), .A2(KEYINPUT35), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(G116), .A3(new_n216), .A4(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n405), .A2(G77), .A3(new_n214), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(G50), .B2(new_n219), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n717), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(G367));
  INV_X1    g0709(.A(KEYINPUT100), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n603), .A2(new_n666), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n709), .A2(new_n711), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n645), .A2(new_n666), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n672), .A2(new_n677), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n617), .B1(new_n912), .B2(new_n591), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n916), .A2(KEYINPUT42), .B1(new_n917), .B2(new_n673), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT99), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT42), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n542), .A2(new_n673), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(new_n552), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n552), .A3(new_n632), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n910), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n922), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n920), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(KEYINPUT100), .A3(new_n932), .A4(new_n918), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n927), .B(KEYINPUT43), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n923), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n676), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(KEYINPUT101), .A3(new_n914), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n914), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT101), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n941), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n682), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n915), .ZN(new_n948));
  INV_X1    g0748(.A(new_n677), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n675), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT106), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n671), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n671), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n950), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT44), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n679), .B2(new_n914), .ZN(new_n958));
  INV_X1    g0758(.A(new_n914), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n678), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT103), .Z(new_n963));
  NAND3_X1  g0763(.A1(new_n679), .A2(new_n914), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n959), .B2(new_n678), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n961), .A2(new_n676), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n955), .A2(new_n956), .A3(new_n715), .A4(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n960), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT44), .B1(new_n959), .B2(new_n678), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n964), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT104), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n961), .A2(KEYINPUT104), .A3(new_n964), .A4(new_n966), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n937), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n676), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n974), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n968), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n715), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n947), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n722), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n945), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n743), .A2(G97), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n746), .A2(G317), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G303), .A2(new_n756), .B1(new_n758), .B2(G283), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n750), .A2(G311), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n760), .A2(new_n459), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n991), .B(new_n274), .C1(new_n580), .C2(new_n770), .ZN(new_n992));
  INV_X1    g0792(.A(new_n764), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n990), .A2(KEYINPUT46), .B1(new_n993), .B2(new_n354), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n989), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT107), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n993), .A2(new_n219), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n274), .B(new_n997), .C1(G143), .C2(new_n750), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G150), .A2(new_n756), .B1(new_n751), .B2(G159), .ZN(new_n999));
  INV_X1    g0799(.A(new_n760), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n252), .A2(new_n1000), .B1(new_n758), .B2(G50), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n597), .A2(new_n742), .B1(new_n745), .B2(new_n797), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n729), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n925), .A2(new_n727), .A3(new_n926), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n238), .A2(new_n732), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n731), .B1(new_n681), .B2(new_n521), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n724), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n984), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(new_n735), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1015), .A2(new_n685), .B1(G107), .B2(new_n210), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n234), .A2(G45), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n361), .A2(new_n202), .ZN(new_n1019));
  XOR2_X1   g0819(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n475), .B1(new_n219), .B2(new_n597), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n681), .B(new_n327), .C1(new_n1024), .C2(new_n685), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1016), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G322), .A2(new_n750), .B1(new_n751), .B2(G311), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n761), .B2(new_n757), .C1(new_n1028), .C2(new_n755), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n993), .A2(new_n792), .B1(new_n760), .B2(new_n580), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT112), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n327), .B1(new_n746), .B2(G326), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n459), .B2(new_n742), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1037), .B2(KEYINPUT49), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n760), .A2(new_n597), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n274), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n985), .B(new_n1043), .C1(new_n798), .C2(new_n745), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT110), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n993), .A2(new_n364), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G68), .A2(new_n758), .B1(new_n750), .B2(G159), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n202), .B2(new_n755), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n253), .C2(new_n751), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1038), .A2(new_n1041), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n723), .B1(new_n731), .B2(new_n1026), .C1(new_n1050), .C2(new_n788), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT113), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n727), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1054), .C1(new_n675), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n955), .A2(new_n956), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n722), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n715), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n955), .A2(new_n715), .A3(new_n956), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n682), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1056), .B(new_n1058), .C1(new_n1059), .C2(new_n1061), .ZN(G393));
  AND2_X1   g0862(.A1(new_n243), .A2(new_n732), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n730), .B1(new_n330), .B2(new_n210), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n723), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n769), .A2(new_n798), .B1(new_n755), .B2(new_n386), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n327), .B1(new_n760), .B2(new_n219), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n770), .A2(new_n202), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n361), .C2(new_n758), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n993), .A2(new_n597), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G87), .A2(new_n743), .B1(new_n746), .B2(G143), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n770), .A2(new_n761), .B1(new_n792), .B2(new_n760), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n327), .B(new_n1075), .C1(G294), .C2(new_n758), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G107), .A2(new_n743), .B1(new_n746), .B2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n459), .C2(new_n993), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n756), .A2(G311), .B1(new_n750), .B2(G317), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1074), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1065), .B1(new_n1081), .B2(new_n729), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n914), .B2(new_n1055), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n971), .A2(new_n937), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n967), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1085), .B2(new_n983), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n968), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n977), .A2(new_n978), .A3(new_n974), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n978), .B1(new_n977), .B2(new_n974), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n683), .B1(new_n1060), .B2(new_n1085), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1089), .A2(new_n1095), .ZN(G390));
  AND2_X1   g0896(.A1(new_n835), .A2(new_n701), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n886), .A2(new_n890), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n892), .A3(new_n893), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n713), .A2(new_n673), .A3(new_n811), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n812), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT116), .B1(new_n1104), .B2(new_n812), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n885), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n890), .B(KEYINPUT115), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n876), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1099), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(new_n812), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n812), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n885), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n876), .A3(new_n1109), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1099), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n1102), .A4(new_n1101), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n983), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT119), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n892), .A2(new_n725), .A3(new_n893), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n786), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n723), .B1(new_n253), .B2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n327), .B(new_n1071), .C1(G87), .C2(new_n1000), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n756), .A2(G116), .B1(new_n750), .B2(G283), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G97), .A2(new_n758), .B1(new_n751), .B2(G107), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G68), .A2(new_n743), .B1(new_n746), .B2(G294), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n769), .A2(new_n1132), .B1(new_n755), .B2(new_n805), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT118), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1000), .A2(G150), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(KEYINPUT53), .B1(G159), .B2(new_n764), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(KEYINPUT53), .C2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n327), .B1(new_n770), .B2(new_n797), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n758), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1141), .B1(new_n202), .B2(new_n742), .C1(new_n1142), .C2(new_n745), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1131), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1144), .B2(new_n729), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1124), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1122), .A2(new_n1123), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT119), .B1(new_n1121), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1098), .B(new_n1097), .C1(new_n1118), .C2(new_n1101), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1119), .A2(new_n1118), .A3(new_n1102), .A4(new_n1101), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n885), .B1(new_n701), .B2(new_n814), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n884), .B1(new_n1097), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n835), .A2(new_n701), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n670), .B(new_n813), .C1(new_n689), .C2(new_n700), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n885), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n456), .A2(new_n701), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n897), .A2(new_n659), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n683), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n1167), .ZN(G378));
  NOR3_X1   g0968(.A1(new_n894), .A2(new_n887), .A3(new_n888), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n877), .A2(new_n876), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n864), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(G330), .C1(new_n862), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n379), .A2(new_n377), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n653), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n268), .A2(new_n838), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT121), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n653), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1177), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT121), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1176), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1174), .A2(new_n1175), .A3(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1172), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n896), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1196), .B2(new_n1173), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n722), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n723), .B1(G50), .B2(new_n1125), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT120), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n274), .A2(new_n287), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n997), .A2(new_n1042), .A3(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n756), .A2(G107), .B1(new_n758), .B2(new_n521), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G116), .A2(new_n750), .B1(new_n751), .B2(G97), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n792), .B2(new_n745), .C1(new_n772), .C2(new_n742), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G50), .B1(new_n254), .B2(new_n287), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1207), .A2(KEYINPUT58), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n769), .A2(new_n1142), .B1(new_n770), .B2(new_n805), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G128), .A2(new_n756), .B1(new_n1000), .B2(new_n1140), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n798), .B2(new_n993), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G137), .C2(new_n758), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n254), .B(new_n287), .C1(new_n742), .C2(new_n386), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G124), .B2(new_n746), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1209), .B1(KEYINPUT58), .B2(new_n1207), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1200), .B1(new_n1220), .B2(new_n729), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1192), .B2(new_n726), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1198), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1192), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1196), .A2(new_n1194), .A3(new_n1173), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1166), .B2(new_n1162), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1163), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1162), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(KEYINPUT122), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1166), .A2(new_n1227), .A3(new_n1162), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT122), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1233), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n683), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1223), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT123), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(KEYINPUT123), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n1160), .A2(new_n722), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n724), .B1(new_n219), .B2(new_n786), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n274), .B1(new_n742), .B2(new_n597), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT125), .Z(new_n1247));
  AOI22_X1  g1047(.A1(G294), .A2(new_n750), .B1(new_n751), .B2(G116), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n792), .B2(new_n755), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n745), .A2(new_n761), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n760), .A2(new_n330), .B1(new_n757), .B2(new_n354), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1249), .A2(new_n1046), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n327), .B1(new_n993), .B2(new_n202), .C1(new_n770), .C2(new_n1139), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n769), .A2(new_n805), .B1(new_n755), .B2(new_n797), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n760), .A2(new_n386), .B1(new_n757), .B2(new_n798), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1132), .A2(new_n745), .B1(new_n742), .B2(new_n772), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1247), .A2(new_n1252), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1245), .B1(new_n788), .B2(new_n1259), .C1(new_n885), .C2(new_n726), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1244), .A2(new_n1260), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n946), .B(KEYINPUT124), .Z(new_n1262));
  AND2_X1   g1062(.A1(new_n1163), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G381));
  NOR4_X1   g1066(.A1(G393), .A2(G390), .A3(G396), .A4(G384), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1013), .A3(new_n1265), .ZN(new_n1268));
  OR3_X1    g1068(.A1(G375), .A2(G378), .A3(new_n1268), .ZN(G407));
  AOI22_X1  g1069(.A1(new_n1147), .A2(new_n1149), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(G343), .C2(new_n1271), .ZN(G409));
  NAND2_X1  g1072(.A1(new_n665), .A2(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1264), .B1(new_n1165), .B2(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1160), .A2(new_n1162), .A3(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n683), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1261), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(G384), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(G384), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1270), .B(new_n1223), .C1(new_n1234), .C2(new_n1239), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1223), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1237), .A2(new_n1226), .A3(new_n1262), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G378), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1273), .B(new_n1281), .C1(new_n1282), .C2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1273), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(G2897), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1281), .B(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1240), .B2(G378), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1289), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1270), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n682), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1226), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1283), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1273), .A4(new_n1281), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1287), .A2(new_n1288), .A3(new_n1294), .A4(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(new_n784), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1087), .A2(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n984), .B2(new_n1012), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n944), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n942), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n936), .B2(new_n938), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n946), .B1(new_n1093), .B2(new_n715), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(new_n722), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n1011), .A3(G390), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1307), .B1(new_n1317), .B2(KEYINPUT127), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  AOI211_X1 g1119(.A(KEYINPUT126), .B(new_n1319), .C1(new_n1309), .C2(new_n1316), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1306), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n984), .A2(new_n1012), .A3(new_n1308), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G390), .B1(new_n1315), .B2(new_n1011), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1317), .A2(new_n1307), .A3(KEYINPUT127), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1305), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1321), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1304), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1330), .B2(new_n1286), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1286), .A2(new_n1330), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1301), .A2(new_n1273), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1292), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1331), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1335), .ZN(G405));
  OR2_X1    g1136(.A1(new_n1240), .A2(new_n1270), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1321), .A2(new_n1327), .A3(new_n1281), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1281), .B1(new_n1321), .B2(new_n1327), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1271), .B(new_n1337), .C1(new_n1338), .C2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1271), .A2(new_n1337), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1281), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1328), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1321), .A2(new_n1327), .A3(new_n1281), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1340), .A2(new_n1345), .ZN(G402));
endmodule


