//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT97), .B(KEYINPUT11), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G1gat), .B2(new_n208), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT98), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT98), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT15), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n221), .A2(KEYINPUT99), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT15), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n214), .B(KEYINPUT100), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n217), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n219), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT101), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(KEYINPUT101), .A3(new_n219), .A4(new_n227), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n232), .A2(new_n233), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n213), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n232), .A2(new_n213), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n232), .B(new_n213), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n238), .B(KEYINPUT13), .Z(new_n244));
  AOI22_X1  g043(.A1(new_n240), .A2(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n207), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n245), .A3(new_n207), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G169gat), .ZN(new_n251));
  INV_X1    g050(.A(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT72), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n253), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(KEYINPUT26), .B2(new_n253), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G183gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n259), .A2(new_n261), .A3(new_n266), .A4(new_n262), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n260), .A2(G183gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n258), .A2(KEYINPUT27), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT70), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n259), .A2(new_n261), .A3(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n272), .A2(KEYINPUT28), .A3(new_n262), .A4(new_n274), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n268), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n269), .B1(new_n268), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n257), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(G127gat), .A2(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G127gat), .A2(G134gat), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT74), .A2(G120gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT74), .A2(G120gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(G113gat), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G120gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n284), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(KEYINPUT73), .A2(G134gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT73), .A2(G134gat), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n279), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n256), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n258), .A2(new_n262), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n301), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT25), .A4(new_n305), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n256), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT24), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n309), .A2(new_n310), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n313), .B1(new_n322), .B2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AOI211_X1 g124(.A(KEYINPUT68), .B(new_n312), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(new_n313), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n312), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n278), .B(new_n299), .C1(new_n326), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n324), .B1(new_n320), .B2(new_n321), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n335), .A2(new_n336), .A3(new_n313), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT68), .B1(new_n337), .B2(new_n312), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n327), .A3(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n299), .B1(new_n340), .B2(new_n278), .ZN(new_n341));
  INV_X1    g140(.A(G227gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n334), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI221_X1 g146(.A(new_n345), .B1(new_n342), .B2(new_n343), .C1(new_n334), .C2(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G71gat), .B(G99gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n278), .B1(new_n326), .B2(new_n332), .ZN(new_n354));
  INV_X1    g153(.A(new_n299), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n342), .A2(new_n343), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n333), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(KEYINPUT76), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n353), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT33), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n350), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n347), .A2(new_n369), .A3(new_n348), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n360), .A2(KEYINPUT76), .A3(new_n361), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT76), .B1(new_n360), .B2(new_n361), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378));
  AND2_X1   g177(.A1(KEYINPUT78), .A2(G211gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT78), .A2(G211gat), .ZN(new_n380));
  OAI21_X1  g179(.A(G218gat), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  OR2_X1    g181(.A1(G197gat), .A2(G204gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(G197gat), .A2(G204gat), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n385), .B2(KEYINPUT79), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT78), .B(G211gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT22), .B1(new_n387), .B2(G218gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n383), .A2(new_n384), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(KEYINPUT79), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G141gat), .B(G148gat), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n398), .B(new_n404), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n396), .B2(new_n405), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n401), .A2(new_n403), .ZN(new_n411));
  AND2_X1   g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n403), .A2(KEYINPUT83), .A3(KEYINPUT2), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n410), .A2(new_n411), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI22_X1  g218(.A1(new_n392), .A2(new_n395), .B1(KEYINPUT29), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n408), .A2(new_n416), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n378), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n394), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n429), .B2(new_n417), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n427), .A2(new_n394), .B1(new_n428), .B2(new_n418), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n422), .B(new_n423), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n417), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n416), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n423), .B1(new_n431), .B2(KEYINPUT88), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n420), .ZN(new_n437));
  AOI21_X1  g236(.A(G22gat), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n377), .B1(new_n438), .B2(KEYINPUT89), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n437), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n437), .A3(G22gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n442), .A2(KEYINPUT89), .A3(new_n443), .A4(new_n377), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n374), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT95), .B1(new_n370), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n349), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT95), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n374), .A4(new_n447), .ZN(new_n453));
  AND2_X1   g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n278), .B(new_n454), .C1(new_n326), .C2(new_n332), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n330), .A2(new_n331), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n278), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n454), .A2(KEYINPUT29), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n392), .A2(new_n395), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n461), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n278), .A2(new_n456), .A3(new_n454), .ZN(new_n464));
  INV_X1    g263(.A(new_n354), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G8gat), .B(G36gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n462), .A2(new_n466), .A3(KEYINPUT30), .A4(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT80), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g278(.A1(G225gat), .A2(G233gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n417), .B1(new_n408), .B2(new_n416), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n419), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n299), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n290), .A2(new_n298), .A3(new_n424), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT86), .B1(new_n485), .B2(KEYINPUT4), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n290), .A2(new_n298), .A3(new_n424), .A4(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT85), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n479), .B(new_n484), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(new_n281), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n284), .A2(new_n287), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n295), .A2(new_n297), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n434), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n485), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n479), .B1(new_n504), .B2(new_n481), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n496), .A2(new_n505), .A3(KEYINPUT84), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT84), .B1(new_n496), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n493), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT0), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G85gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT87), .B(KEYINPUT6), .Z(new_n515));
  OAI211_X1 g314(.A(new_n493), .B(new_n512), .C1(new_n506), .C2(new_n507), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n515), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n462), .A2(new_n466), .A3(new_n470), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT81), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT81), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n462), .A2(new_n466), .A3(new_n524), .A4(new_n470), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n478), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n449), .A2(new_n453), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n369), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n364), .B2(new_n365), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT94), .B(new_n374), .C1(new_n530), .C2(new_n350), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT94), .B1(new_n451), .B2(new_n374), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n445), .A2(new_n446), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n508), .A2(KEYINPUT92), .A3(new_n513), .A4(new_n518), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n472), .A3(new_n473), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n536), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT35), .A2(new_n528), .B1(new_n534), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n503), .A2(new_n480), .A3(new_n485), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(KEYINPUT39), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n494), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n486), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n491), .B(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n550), .A2(new_n552), .B1(new_n299), .B2(new_n483), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n547), .B1(new_n553), .B2(new_n480), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n483), .A2(new_n299), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n489), .B2(new_n492), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT90), .B(KEYINPUT39), .Z(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n481), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT40), .A4(new_n512), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n514), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n552), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n480), .B1(new_n561), .B2(new_n555), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n513), .B1(new_n562), .B2(new_n557), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT40), .B1(new_n563), .B2(new_n554), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n535), .B1(new_n565), .B2(new_n542), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n460), .A2(new_n463), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n461), .B(new_n464), .C1(new_n465), .C2(new_n459), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT37), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n462), .A2(new_n466), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n470), .A2(KEYINPUT38), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT91), .A4(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n522), .A2(new_n525), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n540), .A2(new_n577), .A3(new_n517), .A4(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT38), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n570), .B1(new_n462), .B2(new_n466), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n470), .ZN(new_n582));
  INV_X1    g381(.A(new_n571), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT93), .B1(new_n581), .B2(new_n470), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n566), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n451), .A2(new_n374), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n451), .A2(new_n590), .A3(new_n374), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n478), .A2(new_n520), .A3(new_n526), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n535), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n587), .A2(new_n589), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(new_n545), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n597));
  INV_X1    g396(.A(new_n533), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n544), .A2(new_n598), .A3(new_n531), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n594), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n250), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G57gat), .B(G64gat), .Z(new_n604));
  AND2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n604), .B(KEYINPUT102), .C1(KEYINPUT9), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G71gat), .B(G78gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT104), .B(KEYINPUT19), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n213), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n611), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT20), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT103), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n615), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(G85gat), .ZN(new_n625));
  INV_X1    g424(.A(G92gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(KEYINPUT8), .A2(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT7), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n608), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n612), .A3(new_n635), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n343), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT110), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT110), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n636), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n634), .A2(KEYINPUT106), .A3(new_n635), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT10), .B1(new_n637), .B2(new_n638), .ZN(new_n652));
  OAI22_X1  g451(.A1(new_n651), .A2(new_n652), .B1(new_n640), .B2(new_n343), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n646), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n646), .B2(new_n654), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n650), .B(new_n649), .C1(new_n235), .C2(new_n236), .ZN(new_n663));
  AND3_X1   g462(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n650), .ZN(new_n665));
  INV_X1    g464(.A(new_n232), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n232), .B1(new_n650), .B2(new_n649), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(KEYINPUT107), .A3(new_n664), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n663), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G190gat), .B(G218gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n663), .B(new_n675), .C1(new_n669), .C2(new_n671), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G134gat), .B(G162gat), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n678), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT109), .B(new_n685), .C1(new_n676), .C2(new_n679), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n677), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n236), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n665), .B1(new_n688), .B2(new_n234), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n670), .B2(new_n664), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n668), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT108), .B1(new_n692), .B2(new_n675), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n693), .B2(new_n685), .ZN(new_n694));
  INV_X1    g493(.A(new_n677), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n678), .A3(new_n683), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n623), .B(new_n662), .C1(new_n687), .C2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n603), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n520), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  AND3_X1   g502(.A1(new_n699), .A2(new_n542), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n212), .B1(new_n699), .B2(new_n542), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT42), .B2(new_n704), .ZN(G1325gat));
  INV_X1    g506(.A(G15gat), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n603), .A2(new_n708), .A3(new_n534), .A4(new_n698), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n589), .A2(new_n591), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n699), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n708), .ZN(G1326gat));
  NAND2_X1  g511(.A1(new_n699), .A2(new_n535), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n535), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n718), .B(new_n720), .ZN(G1327gat));
  NAND2_X1  g520(.A1(new_n687), .A2(new_n697), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n596), .B2(new_n602), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n600), .A2(new_n594), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n687), .A2(new_n697), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n623), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n662), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n726), .A2(new_n729), .A3(new_n250), .A4(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n520), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n722), .A2(new_n732), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n603), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n520), .A2(G29gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n738), .A2(new_n736), .A3(new_n739), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(new_n740), .A3(new_n741), .ZN(G1328gat));
  OAI21_X1  g541(.A(G36gat), .B1(new_n734), .B2(new_n543), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n543), .A2(G36gat), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT46), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(G1329gat));
  INV_X1    g546(.A(G43gat), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n603), .A2(new_n748), .A3(new_n534), .A4(new_n737), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n733), .A2(new_n710), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n748), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT47), .B(new_n749), .C1(new_n750), .C2(new_n748), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1330gat));
  NAND2_X1  g554(.A1(new_n535), .A2(G50gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n447), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n734), .A2(new_n756), .B1(new_n757), .B2(G50gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1331gat));
  INV_X1    g559(.A(new_n662), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n728), .A2(new_n249), .A3(new_n623), .A4(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n727), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n700), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n542), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT49), .B(G64gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(G1333gat));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n710), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n532), .A2(new_n533), .A3(G71gat), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n770), .A2(G71gat), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n763), .A2(new_n535), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  OR3_X1    g574(.A1(new_n249), .A2(KEYINPUT114), .A3(new_n730), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT114), .B1(new_n249), .B2(new_n730), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n662), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n726), .A2(new_n729), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n700), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n728), .B(new_n778), .C1(new_n545), .C2(new_n595), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n728), .A4(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n662), .A2(new_n700), .A3(new_n625), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n781), .A2(new_n625), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n761), .A2(G92gat), .A3(new_n543), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n784), .B2(new_n785), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n726), .A2(new_n729), .A3(new_n543), .A4(new_n779), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n790), .B(new_n794), .C1(new_n795), .C2(new_n626), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT115), .B(new_n794), .C1(new_n795), .C2(new_n626), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n545), .A2(new_n595), .A3(KEYINPUT96), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n601), .B1(new_n600), .B2(new_n594), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n724), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n727), .A2(new_n728), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n723), .ZN(new_n806));
  INV_X1    g605(.A(new_n779), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n804), .A2(new_n806), .A3(new_n542), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n793), .B1(new_n808), .B2(G92gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT115), .B1(new_n809), .B2(new_n790), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n799), .B1(new_n801), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(G1337gat));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n786), .A2(new_n813), .A3(new_n534), .A4(new_n662), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n780), .A2(new_n710), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1338gat));
  INV_X1    g615(.A(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n662), .A2(new_n535), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n787), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n780), .A2(G106gat), .A3(new_n535), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1339gat));
  NOR2_X1   g624(.A1(new_n651), .A2(new_n652), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n641), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n653), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n653), .A2(KEYINPUT54), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n658), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n659), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT55), .A4(new_n658), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n238), .B1(new_n237), .B2(new_n239), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n243), .A2(new_n244), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n206), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n832), .A2(new_n248), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n687), .A2(new_n697), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n623), .ZN(new_n839));
  INV_X1    g638(.A(new_n248), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n833), .B(new_n832), .C1(new_n840), .C2(new_n246), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n662), .A2(new_n248), .A3(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n722), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n839), .A2(new_n843), .B1(new_n698), .B2(new_n250), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n844), .B2(new_n535), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n722), .A2(new_n250), .A3(new_n730), .A4(new_n761), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n722), .A2(new_n841), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n623), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n447), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n845), .A2(new_n534), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n542), .A2(new_n520), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n286), .A3(new_n250), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n449), .A2(new_n849), .A3(new_n453), .A4(new_n853), .ZN(new_n856));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n249), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(G1340gat));
  OAI21_X1  g657(.A(G120gat), .B1(new_n854), .B2(new_n761), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n856), .A2(new_n282), .A3(new_n283), .A4(new_n662), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n854), .B2(new_n623), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n856), .A2(new_n294), .A3(new_n730), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1342gat));
  NAND2_X1  g663(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n856), .A2(new_n293), .A3(new_n728), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n854), .B2(new_n722), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1343gat));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  INV_X1    g670(.A(new_n853), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n710), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n250), .A2(G141gat), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n849), .A2(new_n535), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n873), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n447), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n843), .A2(KEYINPUT120), .A3(new_n623), .A4(new_n838), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n846), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n839), .B2(new_n843), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n877), .B1(new_n844), .B2(new_n447), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n250), .B(new_n876), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G141gat), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n871), .B(new_n875), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n875), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT122), .A3(KEYINPUT58), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT122), .B1(new_n889), .B2(KEYINPUT58), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(G1344gat));
  NOR3_X1   g691(.A1(new_n844), .A2(new_n447), .A3(new_n876), .ZN(new_n893));
  INV_X1    g692(.A(G148gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n662), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n882), .A2(new_n883), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n873), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n761), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n894), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n844), .A2(new_n447), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n883), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n662), .A3(new_n873), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n900), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n899), .B2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n897), .B2(new_n623), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n893), .A2(new_n399), .A3(new_n730), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n400), .A3(new_n728), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  OAI21_X1  g710(.A(G162gat), .B1(new_n897), .B2(new_n722), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n543), .A2(new_n700), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n845), .A2(new_n534), .A3(new_n851), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n250), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n449), .A2(new_n453), .A3(new_n542), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR4_X1   g719(.A1(new_n844), .A2(new_n700), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n251), .A3(new_n249), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT125), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n915), .B2(new_n761), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n252), .A3(new_n662), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  NOR2_X1   g726(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n915), .B2(new_n623), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n921), .A2(new_n272), .A3(new_n274), .A4(new_n730), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n921), .A2(new_n262), .A3(new_n728), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n852), .A2(new_n728), .A3(new_n914), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n710), .A2(new_n700), .A3(new_n543), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n901), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n249), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n903), .A2(new_n940), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n249), .A2(G197gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  AOI21_X1  g746(.A(G204gat), .B1(new_n947), .B2(KEYINPUT62), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n662), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n949), .B(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n943), .B2(new_n761), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1353gat));
  NOR2_X1   g752(.A1(new_n623), .A2(new_n387), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n941), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n903), .A2(new_n730), .A3(new_n940), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n943), .B2(new_n722), .ZN(new_n960));
  INV_X1    g759(.A(G218gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n961), .A3(new_n728), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1355gat));
endmodule


