//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT75), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(new_n190), .A3(new_n193), .A4(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(new_n188), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(G146), .A3(new_n194), .A4(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT74), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT68), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G119), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n212), .A2(G119), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n209), .A2(new_n210), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT23), .B1(new_n212), .B2(G119), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n216), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .A4(new_n214), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(new_n203), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n198), .B(new_n202), .C1(new_n218), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT74), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT74), .B1(new_n204), .B2(new_n206), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT68), .A2(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT68), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n216), .B1(new_n231), .B2(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(new_n221), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n228), .A2(new_n232), .B1(new_n233), .B2(G110), .ZN(new_n234));
  INV_X1    g048(.A(new_n198), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n191), .A2(KEYINPUT75), .B1(new_n196), .B2(new_n195), .ZN(new_n236));
  AOI21_X1  g050(.A(G146), .B1(new_n236), .B2(new_n194), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n228), .A2(new_n232), .B1(new_n233), .B2(G110), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n202), .A4(new_n198), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n225), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n243), .A2(KEYINPUT22), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(KEYINPUT22), .ZN(new_n245));
  AOI21_X1  g059(.A(G137), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(G137), .A3(new_n245), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G902), .ZN(new_n251));
  INV_X1    g065(.A(new_n248), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(new_n246), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n225), .A2(new_n238), .A3(new_n240), .A4(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT25), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n250), .A2(new_n257), .A3(new_n251), .A4(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(G217), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(G234), .B2(new_n251), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(G902), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n254), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT77), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(KEYINPUT77), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  AOI21_X1  g084(.A(G131), .B1(new_n269), .B2(G137), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n271), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n200), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(G143), .B2(new_n200), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n231), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n280), .B2(G146), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n200), .A2(KEYINPUT66), .A3(G143), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n281), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G131), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n272), .A2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n269), .A2(G137), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n278), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT0), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n212), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n299), .A2(new_n212), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n304), .A3(new_n282), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n287), .A2(new_n303), .A3(new_n281), .A4(new_n288), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n270), .A2(new_n273), .A3(new_n294), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n278), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n267), .B1(new_n297), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n278), .A2(new_n309), .ZN(new_n312));
  INV_X1    g126(.A(new_n307), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n295), .B1(new_n275), .B2(new_n277), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n213), .A2(new_n214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n279), .A2(KEYINPUT1), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n317), .A2(new_n318), .B1(new_n279), .B2(new_n281), .ZN(new_n319));
  AND4_X1   g133(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n281), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n290), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n314), .A2(new_n323), .A3(KEYINPUT30), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g139(.A1(G116), .A2(G119), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(G116), .A2(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G116), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT69), .A3(new_n326), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT2), .B(G113), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n326), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n311), .A2(new_n324), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(KEYINPUT71), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n314), .A2(new_n323), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT26), .B(G101), .ZN(new_n345));
  NOR2_X1   g159(.A1(G237), .A2(G953), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G210), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT31), .B1(new_n340), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n339), .B1(new_n297), .B2(new_n310), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n290), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT70), .B1(new_n285), .B2(new_n290), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n310), .B1(new_n359), .B2(new_n315), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n343), .A2(new_n342), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT28), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n350), .B1(new_n356), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n350), .B1(new_n360), .B2(new_n362), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n311), .A2(new_n324), .A3(new_n339), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n353), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n370), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n351), .B1(new_n356), .B2(new_n363), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(new_n344), .A3(new_n350), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n344), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n314), .A2(new_n323), .B1(new_n342), .B2(new_n343), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n363), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n251), .ZN(new_n384));
  OAI21_X1  g198(.A(G472), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n373), .A2(new_n374), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n373), .A2(new_n385), .A3(KEYINPUT73), .A4(new_n374), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n266), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n199), .A2(new_n200), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n201), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n242), .A3(G214), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n280), .ZN(new_n395));
  NAND2_X1  g209(.A1(G143), .A2(G214), .ZN(new_n396));
  NOR4_X1   g210(.A1(new_n396), .A2(KEYINPUT85), .A3(G237), .A4(G953), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n398));
  AND2_X1   g212(.A1(G143), .A2(G214), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n346), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n395), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n242), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT85), .B1(new_n405), .B2(new_n396), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n346), .A3(new_n398), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n395), .A3(new_n402), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n392), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n192), .A2(new_n194), .A3(new_n197), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n200), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(KEYINPUT17), .A3(G131), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(new_n198), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(G131), .B1(new_n394), .B2(new_n280), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n400), .B2(new_n397), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT86), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n401), .A2(G131), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n420), .A3(new_n415), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n410), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(G104), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT87), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n392), .A2(new_n404), .A3(new_n409), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT19), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n199), .B(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n198), .B1(new_n430), .B2(G146), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n423), .A2(new_n426), .B1(new_n432), .B2(new_n425), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT20), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n422), .A2(new_n198), .A3(new_n412), .A4(new_n413), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n427), .A3(new_n426), .ZN(new_n438));
  AOI22_X1  g252(.A1(KEYINPUT86), .A2(new_n416), .B1(new_n401), .B2(G131), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n431), .B1(new_n421), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n425), .B1(new_n440), .B2(new_n410), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n434), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n437), .A2(new_n427), .A3(new_n426), .ZN(new_n446));
  INV_X1    g260(.A(new_n425), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n437), .B2(new_n427), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n251), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G475), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n213), .A2(G143), .A3(new_n214), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n280), .A2(G128), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n454), .A2(G134), .B1(new_n455), .B2(new_n452), .ZN(new_n456));
  AND4_X1   g270(.A1(KEYINPUT13), .A2(new_n452), .A3(G134), .A4(new_n455), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT88), .B1(new_n330), .B2(G122), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n330), .A2(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G107), .ZN(new_n465));
  INV_X1    g279(.A(G107), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n456), .A2(new_n457), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n469), .A3(G107), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n462), .B(new_n463), .C1(KEYINPUT14), .C2(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n455), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n269), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n452), .A2(G134), .A3(new_n455), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n470), .A2(new_n471), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n476), .A2(new_n259), .A3(G953), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n468), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n468), .B2(new_n475), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n251), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT89), .B(new_n251), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n486), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(G234), .A2(G237), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n491), .A2(G952), .A3(new_n242), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n491), .A2(G902), .A3(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n451), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n466), .A2(G104), .ZN(new_n498));
  AND2_X1   g312(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n499));
  NOR2_X1   g313(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(G104), .A3(new_n466), .ZN(new_n504));
  INV_X1    g318(.A(G104), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G107), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n466), .A2(G104), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n505), .A2(G107), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n503), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n502), .B1(new_n511), .B2(new_n501), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n514));
  INV_X1    g328(.A(new_n501), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n504), .A2(new_n506), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(G101), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n339), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT82), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G101), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n339), .A4(new_n517), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT5), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n331), .A3(G116), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n329), .A2(new_n333), .ZN(new_n526));
  OAI211_X1 g340(.A(G113), .B(new_n525), .C1(new_n526), .C2(new_n524), .ZN(new_n527));
  OAI21_X1  g341(.A(G101), .B1(new_n510), .B2(new_n509), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n507), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n338), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n519), .A2(new_n530), .A3(new_n532), .A4(new_n523), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT6), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT84), .B1(new_n313), .B2(new_n189), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n319), .A2(new_n320), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n189), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n313), .A2(KEYINPUT84), .A3(new_n189), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n544), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n534), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n535), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n534), .A2(KEYINPUT6), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n538), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n542), .B2(new_n543), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n507), .A2(new_n528), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n527), .A2(new_n338), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n525), .A2(G113), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n524), .B1(new_n332), .B2(new_n326), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n338), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n529), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n532), .B(KEYINPUT8), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n542), .A2(new_n543), .A3(new_n552), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n564), .B2(new_n535), .ZN(new_n565));
  OAI21_X1  g379(.A(G210), .B1(G237), .B2(G902), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n551), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n551), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n497), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n242), .A2(G227), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G140), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT78), .B(G110), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n287), .A2(new_n281), .A3(new_n288), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n318), .A2(G128), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n320), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(new_n554), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n578), .A2(new_n577), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n507), .B(new_n528), .C1(new_n583), .C2(new_n320), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT80), .A3(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n312), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n554), .A2(new_n576), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n307), .B1(new_n514), .B2(new_n512), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n359), .A2(new_n588), .B1(new_n589), .B2(new_n521), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT81), .B1(new_n529), .B2(new_n291), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT81), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n540), .A2(new_n554), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n584), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n595), .A2(KEYINPUT12), .A3(new_n312), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT12), .B1(new_n595), .B2(new_n312), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n575), .B(new_n591), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n586), .A2(new_n590), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n312), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n575), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n570), .B(new_n251), .C1(new_n599), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n575), .A3(new_n591), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n586), .A2(new_n590), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n595), .A2(new_n312), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(KEYINPUT12), .A3(new_n312), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n587), .A2(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(G469), .B(new_n604), .C1(new_n610), .C2(new_n575), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n570), .A2(new_n251), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(G221), .B1(new_n476), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n569), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n390), .A2(new_n496), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(new_n451), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n478), .B2(new_n479), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n468), .A2(new_n475), .ZN(new_n623));
  INV_X1    g437(.A(new_n477), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n468), .A2(new_n477), .A3(new_n475), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(KEYINPUT33), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n627), .A3(G478), .A4(new_n251), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n480), .A2(new_n485), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(KEYINPUT90), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT90), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n495), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n569), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n369), .A2(new_n251), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n371), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n616), .A2(new_n266), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT91), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n497), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n551), .A2(new_n565), .ZN(new_n646));
  INV_X1    g460(.A(new_n566), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n551), .A2(new_n565), .A3(new_n566), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT93), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n436), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT92), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n653), .B(KEYINPUT20), .C1(new_n433), .C2(new_n435), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n486), .B1(new_n482), .B2(new_n483), .ZN(new_n656));
  INV_X1    g470(.A(new_n489), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n450), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n650), .A2(new_n651), .A3(new_n634), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n634), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT93), .B1(new_n569), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n640), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n253), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT94), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n253), .A2(new_n667), .A3(new_n668), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n249), .A2(KEYINPUT95), .A3(KEYINPUT36), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT94), .B1(new_n674), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n241), .ZN(new_n677));
  INV_X1    g491(.A(new_n241), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n262), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n261), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n496), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n639), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n617), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT37), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT96), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G110), .ZN(G12));
  NAND2_X1  g501(.A1(new_n388), .A2(new_n389), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n614), .A2(new_n615), .A3(new_n681), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n492), .B1(new_n493), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n659), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n688), .A2(new_n694), .A3(new_n650), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT97), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n655), .A2(new_n658), .A3(new_n691), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n615), .A3(new_n614), .A4(new_n681), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n569), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT97), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n688), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  INV_X1    g517(.A(new_n616), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n691), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n648), .A2(new_n649), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT38), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n378), .A2(new_n351), .A3(new_n379), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(G902), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n350), .B1(new_n366), .B2(new_n344), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n373), .A2(new_n374), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT98), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n373), .A2(new_n716), .A3(new_n713), .A4(new_n374), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n490), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n620), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n497), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n718), .A2(new_n681), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n707), .A2(new_n709), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n280), .ZN(G45));
  AOI21_X1  g539(.A(new_n689), .B1(new_n388), .B2(new_n389), .ZN(new_n726));
  INV_X1    g540(.A(new_n632), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n451), .A3(new_n692), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n569), .A2(new_n728), .A3(KEYINPUT100), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT100), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n620), .A2(new_n632), .A3(new_n691), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n730), .B1(new_n650), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n726), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NOR2_X1   g548(.A1(new_n570), .A2(KEYINPUT101), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n599), .A2(new_n602), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n736), .B2(G902), .ZN(new_n737));
  OAI221_X1 g551(.A(new_n251), .B1(KEYINPUT101), .B2(new_n570), .C1(new_n599), .C2(new_n602), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n615), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n390), .A2(new_n636), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  INV_X1    g557(.A(new_n266), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n370), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT32), .B1(new_n369), .B2(new_n370), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT73), .B1(new_n747), .B2(new_n385), .ZN(new_n748));
  INV_X1    g562(.A(new_n389), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n744), .B(new_n740), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n660), .B2(new_n662), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT102), .B(G116), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G18));
  AOI21_X1  g567(.A(new_n682), .B1(new_n388), .B2(new_n389), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n569), .A2(new_n739), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  OAI211_X1 g571(.A(new_n720), .B(new_n497), .C1(new_n567), .C2(new_n568), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n370), .B(KEYINPUT103), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n353), .A2(new_n368), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n351), .B1(new_n380), .B2(new_n381), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n744), .A2(new_n638), .A3(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n739), .A3(new_n495), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  AND3_X1   g581(.A1(new_n365), .A2(new_n367), .A3(new_n366), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n367), .B1(new_n365), .B2(new_n366), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(G902), .B1(new_n770), .B2(new_n364), .ZN(new_n771));
  INV_X1    g585(.A(G472), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n681), .B(new_n763), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n638), .A2(KEYINPUT104), .A3(new_n681), .A4(new_n763), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n728), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n755), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n189), .ZN(G27));
  NOR3_X1   g593(.A1(new_n708), .A2(new_n616), .A3(new_n645), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n390), .A2(new_n780), .A3(new_n731), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n266), .B1(new_n747), .B2(new_n385), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n731), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n781), .A2(new_n782), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n292), .ZN(G33));
  XNOR2_X1  g600(.A(new_n693), .B(KEYINPUT106), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n390), .A3(new_n780), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  NAND2_X1  g603(.A1(new_n727), .A2(new_n620), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n639), .A2(new_n681), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT44), .Z(new_n794));
  OR2_X1    g608(.A1(new_n610), .A2(new_n575), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n604), .ZN(new_n796));
  OAI21_X1  g610(.A(G469), .B1(new_n796), .B2(KEYINPUT45), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n795), .A2(KEYINPUT45), .A3(new_n604), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n613), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT46), .B(new_n613), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n603), .A3(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n803), .A2(new_n615), .A3(new_n705), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n708), .A2(new_n645), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT107), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n803), .A2(new_n810), .A3(new_n615), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n803), .B2(new_n615), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n811), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n688), .A2(new_n744), .A3(new_n728), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n805), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NAND2_X1  g634(.A1(new_n737), .A2(new_n738), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT49), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n615), .A2(new_n497), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n822), .A2(new_n266), .A3(new_n790), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n709), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n718), .ZN(new_n826));
  INV_X1    g640(.A(G952), .ZN(new_n827));
  INV_X1    g641(.A(new_n492), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n791), .A2(new_n828), .A3(new_n764), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n827), .B(G953), .C1(new_n829), .C2(new_n755), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n791), .A2(new_n828), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n805), .A2(new_n740), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n783), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n830), .B(new_n836), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n718), .A2(new_n744), .A3(new_n492), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n832), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n839), .B2(new_n832), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n633), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n620), .A3(new_n632), .A4(new_n841), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n775), .A2(new_n776), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n831), .A2(new_n845), .A3(new_n833), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n645), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n739), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n829), .A2(new_n825), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n844), .B(new_n846), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n821), .A2(new_n615), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n814), .A2(new_n816), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n829), .A2(new_n806), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n843), .B1(new_n857), .B2(KEYINPUT51), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n859), .B(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n261), .A2(new_n680), .A3(new_n692), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n614), .A2(new_n615), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n715), .B2(new_n717), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n759), .A2(new_n864), .B1(new_n777), .B2(new_n755), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n700), .A2(new_n688), .A3(new_n694), .A4(new_n650), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n700), .B1(new_n699), .B2(new_n688), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n733), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n702), .A2(KEYINPUT111), .A3(new_n733), .A4(new_n865), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n663), .A2(new_n390), .A3(new_n740), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n755), .A2(new_n754), .B1(new_n759), .B2(new_n765), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n741), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n719), .A2(new_n451), .A3(new_n495), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n650), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT110), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT110), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n650), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n640), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n633), .B(KEYINPUT109), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n640), .A3(new_n634), .A4(new_n650), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n618), .A3(new_n684), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n450), .A2(new_n692), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n655), .A2(new_n490), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n726), .A2(new_n805), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n780), .A2(new_n777), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n788), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n785), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n877), .A2(new_n878), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n891), .A2(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n874), .A2(new_n869), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n872), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n899), .B(KEYINPUT54), .C1(new_n878), .C2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n890), .A2(new_n896), .A3(new_n878), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n741), .A2(new_n756), .A3(new_n766), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT113), .B1(new_n906), .B2(new_n751), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT113), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n879), .A2(new_n880), .A3(new_n908), .A4(new_n741), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n785), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g726(.A(KEYINPUT114), .B(new_n785), .C1(new_n907), .C2(new_n909), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n872), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT52), .B1(new_n872), .B2(new_n873), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n898), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n914), .A2(new_n877), .B1(new_n917), .B2(new_n878), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n861), .A2(new_n904), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n827), .A2(new_n242), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n921), .A2(new_n922), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n826), .B1(new_n925), .B2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n918), .A2(new_n251), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G210), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n538), .A2(new_n549), .A3(new_n550), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n548), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT119), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n242), .A2(G952), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G51));
  NAND2_X1  g753(.A1(new_n914), .A2(new_n877), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n917), .A2(new_n878), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT54), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n918), .A2(new_n919), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n612), .B(KEYINPUT57), .Z(new_n946));
  OAI22_X1  g760(.A1(new_n945), .A2(new_n946), .B1(new_n602), .B2(new_n599), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n797), .A2(new_n798), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n928), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n938), .B1(new_n947), .B2(new_n949), .ZN(G54));
  NAND3_X1  g764(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n951), .A2(new_n433), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n433), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n938), .ZN(G60));
  NAND2_X1  g768(.A1(new_n622), .A2(new_n627), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n943), .B2(new_n944), .ZN(new_n959));
  INV_X1    g773(.A(new_n938), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(KEYINPUT121), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  INV_X1    g776(.A(new_n958), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n942), .A2(KEYINPUT54), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n920), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n965), .B2(new_n938), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n920), .A2(new_n904), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n955), .B1(new_n967), .B2(new_n957), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n961), .A2(new_n966), .A3(new_n968), .ZN(G63));
  XNOR2_X1  g783(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT123), .B1(new_n918), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n250), .A2(new_n254), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  INV_X1    g789(.A(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n903), .A2(KEYINPUT53), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n876), .A2(new_n912), .A3(new_n913), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n973), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n960), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n677), .A2(new_n679), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n973), .B2(new_n979), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n970), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n973), .A2(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n982), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(KEYINPUT61), .A3(new_n960), .A4(new_n980), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n984), .A2(new_n988), .ZN(G66));
  NOR3_X1   g803(.A1(new_n494), .A2(new_n545), .A3(new_n242), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n891), .B2(new_n242), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n930), .B1(G898), .B2(new_n242), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n804), .A2(new_n759), .A3(new_n783), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n807), .A2(new_n995), .A3(new_n788), .ZN(new_n996));
  INV_X1    g810(.A(new_n702), .ZN(new_n997));
  INV_X1    g811(.A(new_n733), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n997), .A2(new_n998), .A3(new_n778), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n996), .A2(new_n785), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n819), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n311), .A2(new_n324), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(new_n430), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n690), .A2(KEYINPUT125), .A3(G227), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT125), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n1006), .B2(G900), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1004), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n888), .B1(new_n620), .B2(new_n490), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(new_n706), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n390), .A3(new_n805), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n807), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OR3_X1    g831(.A1(new_n724), .A2(KEYINPUT62), .A3(new_n999), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT62), .B1(new_n724), .B2(new_n999), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1017), .A2(new_n819), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n994), .B(new_n1010), .C1(new_n1022), .C2(new_n1004), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1004), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g838(.A(KEYINPUT126), .B1(new_n1024), .B2(new_n1009), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(G72));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  NAND2_X1  g842(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n891), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1018), .A2(new_n819), .A3(new_n1019), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n712), .ZN(new_n1033));
  INV_X1    g847(.A(new_n376), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1028), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1034), .A2(new_n712), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT127), .Z(new_n1037));
  OAI211_X1 g851(.A(new_n899), .B(new_n1037), .C1(new_n878), .C2(new_n903), .ZN(new_n1038));
  INV_X1    g852(.A(new_n891), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1028), .B1(new_n1001), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n938), .B1(new_n1040), .B2(new_n1034), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1033), .A2(new_n1038), .A3(new_n1041), .ZN(G57));
endmodule


