//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT85), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT75), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n213), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n207), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n214), .A2(new_n217), .B1(new_n207), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n206), .B1(new_n218), .B2(KEYINPUT29), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G162gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT78), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G141gat), .B(G148gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT79), .B(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n227), .B2(new_n222), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT78), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n223), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n214), .A2(new_n217), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT74), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n209), .A2(new_n240), .A3(new_n213), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n207), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G228gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT86), .B(G22gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT29), .B1(new_n238), .B2(new_n242), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n234), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g050(.A(new_n247), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n248), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n249), .B1(new_n248), .B2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n205), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n253), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(G22gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n258), .B2(G22gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n248), .A2(KEYINPUT88), .A3(new_n249), .A4(new_n253), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n204), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n257), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT0), .ZN(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  INV_X1    g074(.A(G134gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G127gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  INV_X1    g078(.A(G120gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G113gat), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G120gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT70), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285));
  OR3_X1    g084(.A1(new_n280), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n279), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n277), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n281), .A2(new_n283), .ZN(new_n292));
  OAI221_X1 g091(.A(new_n291), .B1(new_n290), .B2(new_n275), .C1(new_n292), .C2(KEYINPUT1), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n289), .A2(new_n233), .A3(new_n230), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT4), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT78), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n297), .A2(new_n224), .A3(new_n225), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n298), .A2(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n293), .A4(new_n289), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n299), .A2(new_n206), .B1(new_n293), .B2(new_n289), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT80), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT80), .B(new_n206), .C1(new_n230), .C2(new_n233), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n294), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n302), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n279), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n284), .A2(new_n286), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n286), .A3(new_n285), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n293), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n234), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(new_n294), .A3(KEYINPUT82), .ZN(new_n318));
  INV_X1    g117(.A(new_n308), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n289), .A2(new_n293), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n234), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n310), .A2(KEYINPUT5), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n307), .A2(new_n325), .A3(new_n308), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n295), .A2(new_n327), .A3(new_n301), .ZN(new_n328));
  INV_X1    g127(.A(new_n320), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(KEYINPUT83), .A3(new_n300), .A4(new_n299), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT6), .B(new_n273), .C1(new_n324), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n336), .B2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(KEYINPUT28), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT26), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n342), .A2(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G226gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G169gat), .ZN(new_n353));
  INV_X1    g152(.A(G176gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT23), .ZN(new_n355));
  AND3_X1   g154(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT66), .B1(new_n341), .B2(KEYINPUT23), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n360), .B(new_n361), .C1(G169gat), .C2(G176gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G190gat), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n338), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n366));
  OR2_X1    g165(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n363), .B(new_n368), .C1(KEYINPUT65), .C2(KEYINPUT25), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n359), .A2(new_n362), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n345), .A2(new_n346), .B1(KEYINPUT23), .B2(new_n341), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT65), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n369), .A2(KEYINPUT68), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT68), .B1(new_n369), .B2(new_n375), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n349), .B(new_n352), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n375), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n374), .B2(new_n373), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n349), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n243), .ZN(new_n385));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT76), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT77), .Z(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n352), .ZN(new_n392));
  AOI221_X4 g191(.A(new_n392), .B1(new_n340), .B2(new_n348), .C1(new_n369), .C2(new_n375), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n349), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n379), .B2(new_n380), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n369), .A2(KEYINPUT68), .A3(new_n375), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n382), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n394), .B(new_n244), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n391), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n310), .B1(new_n326), .B2(new_n331), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n272), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n310), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n326), .A2(new_n331), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n407), .A2(new_n272), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n333), .B(new_n402), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n349), .B1(new_n376), .B2(new_n377), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n393), .B1(new_n413), .B2(new_n382), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n414), .B2(new_n243), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n384), .A2(new_n244), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT91), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n385), .A2(new_n401), .A3(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT38), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n390), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n412), .B1(new_n385), .B2(new_n401), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n390), .A3(new_n422), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n421), .A2(new_n425), .B1(new_n428), .B2(KEYINPUT38), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n268), .B1(new_n411), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n243), .B(new_n393), .C1(new_n413), .C2(new_n382), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n244), .B1(new_n378), .B2(new_n383), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n390), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n402), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n385), .A2(new_n391), .A3(new_n435), .A4(new_n401), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n434), .A2(KEYINPUT89), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT89), .B1(new_n434), .B2(new_n436), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT40), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n319), .B1(new_n318), .B2(new_n322), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n328), .A2(new_n307), .A3(new_n330), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n319), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n441), .A3(new_n319), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n272), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n273), .B1(new_n324), .B2(new_n332), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n443), .A2(new_n319), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n442), .A2(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n440), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n272), .A3(new_n452), .A4(new_n445), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n437), .A2(new_n438), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n413), .A2(new_n329), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n320), .B(new_n349), .C1(new_n376), .C2(new_n377), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT64), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n461), .B(KEYINPUT32), .C1(new_n463), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n457), .A2(new_n458), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT72), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n399), .A2(new_n320), .ZN(new_n476));
  INV_X1    g275(.A(new_n458), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT34), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n472), .A2(new_n480), .A3(new_n473), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(KEYINPUT72), .A2(new_n474), .B1(new_n478), .B2(KEYINPUT34), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(new_n468), .A3(new_n470), .A4(new_n481), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(KEYINPUT73), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  INV_X1    g286(.A(new_n482), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n468), .A4(new_n470), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n483), .A2(KEYINPUT36), .A3(new_n485), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT84), .B1(new_n406), .B2(new_n409), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n405), .A2(new_n272), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n448), .A2(new_n495), .A3(new_n496), .A4(new_n403), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n497), .A3(new_n333), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n434), .A2(new_n436), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n268), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n456), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n490), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n437), .A2(new_n438), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n333), .B1(new_n406), .B2(new_n409), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n267), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n267), .A2(new_n485), .ZN(new_n510));
  INV_X1    g309(.A(new_n483), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(new_n499), .ZN(new_n513));
  INV_X1    g312(.A(new_n333), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n448), .A2(new_n495), .A3(new_n403), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(KEYINPUT84), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n516), .B2(new_n497), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G57gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G64gat), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(G64gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT9), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G71gat), .ZN(new_n524));
  INV_X1    g323(.A(G78gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(KEYINPUT9), .B2(new_n527), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT95), .B(G57gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n521), .B1(new_n532), .B2(G64gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n533), .B2(KEYINPUT96), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(KEYINPUT96), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n529), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT20), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n543), .ZN(new_n545));
  XOR2_X1   g344(.A(G183gat), .B(G211gat), .Z(new_n546));
  OR3_X1    g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G1gat), .B2(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n537), .B2(new_n538), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n547), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n547), .B2(new_n557), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT14), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n567), .A2(KEYINPUT93), .B1(new_n562), .B2(new_n563), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n567), .A2(KEYINPUT93), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT15), .B(new_n561), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n561), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT94), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(KEYINPUT17), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  INV_X1    g381(.A(G99gat), .ZN(new_n583));
  INV_X1    g382(.A(G106gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT8), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT99), .B(G85gat), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n582), .B(new_n585), .C1(G92gat), .C2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n579), .A2(new_n580), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT98), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT41), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n587), .A2(new_n588), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n587), .A2(new_n588), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n597), .B2(new_n577), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n590), .A2(new_n603), .A3(new_n598), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n590), .A2(KEYINPUT100), .A3(new_n603), .A4(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(KEYINPUT101), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n276), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G162gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n605), .A2(new_n608), .A3(new_n612), .A4(new_n606), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n560), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n579), .A2(new_n553), .A3(new_n580), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n553), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n577), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n619), .A2(new_n622), .A3(KEYINPUT18), .A4(new_n620), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n620), .B(KEYINPUT13), .Z(new_n627));
  INV_X1    g426(.A(new_n622), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n621), .A2(new_n577), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT92), .B(G197gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT11), .B(G169gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n625), .A2(new_n630), .A3(new_n626), .A4(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n589), .A2(new_n537), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n589), .A2(new_n537), .ZN(new_n648));
  OAI211_X1 g447(.A(KEYINPUT102), .B(KEYINPUT10), .C1(new_n589), .C2(new_n537), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n647), .ZN(new_n651));
  INV_X1    g450(.A(new_n648), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n644), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n650), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n650), .B2(new_n653), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n618), .A2(new_n642), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n519), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n498), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n663), .A2(new_n504), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n552), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n667), .A2(new_n552), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n491), .B2(new_n492), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n491), .A2(new_n674), .A3(new_n492), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n663), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n503), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n677), .A2(G15gat), .B1(new_n663), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT105), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n268), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  NOR3_X1   g483(.A1(new_n560), .A2(new_n642), .A3(new_n661), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n519), .A2(new_n616), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n562), .A3(new_n664), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n456), .A2(new_n493), .A3(new_n501), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n267), .B(new_n506), .C1(new_n437), .C2(new_n438), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n490), .B2(new_n486), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n518), .B1(new_n692), .B2(KEYINPUT35), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n616), .C1(new_n690), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n493), .A2(KEYINPUT104), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n430), .A2(new_n455), .B1(new_n500), .B2(new_n268), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n491), .A2(new_n674), .A3(new_n492), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n507), .A2(new_n508), .B1(new_n517), .B2(new_n512), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n617), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n694), .B(new_n685), .C1(new_n700), .C2(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n498), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n689), .A2(new_n702), .ZN(G1328gat));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n563), .A3(new_n504), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT46), .Z(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n701), .B2(new_n505), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  NOR2_X1   g506(.A1(new_n676), .A2(new_n675), .ZN(new_n708));
  OAI21_X1  g507(.A(G43gat), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n678), .A2(G43gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n519), .A2(new_n616), .A3(new_n685), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT108), .B(KEYINPUT47), .C1(new_n709), .C2(new_n714), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(G1330gat));
  AND2_X1   g518(.A1(new_n686), .A2(new_n268), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n268), .A2(G50gat), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n720), .A2(G50gat), .B1(new_n701), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g522(.A1(new_n642), .A2(new_n661), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n618), .B(new_n724), .C1(new_n698), .C2(new_n699), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n664), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(new_n532), .Z(G1332gat));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n504), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT49), .B(G64gat), .Z(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1333gat));
  XNOR2_X1  g530(.A(new_n503), .B(KEYINPUT109), .ZN(new_n732));
  AOI21_X1  g531(.A(G71gat), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n708), .A2(new_n524), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n725), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n268), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g537(.A1(new_n560), .A2(new_n641), .A3(new_n660), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n694), .B(new_n739), .C1(new_n700), .C2(KEYINPUT44), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n586), .B1(new_n740), .B2(new_n498), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n560), .A2(new_n641), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n422), .A2(new_n390), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT38), .B1(new_n743), .B2(new_n426), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n419), .B1(new_n415), .B2(new_n416), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n394), .B(new_n243), .C1(new_n399), .C2(new_n400), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n419), .A2(new_n416), .A3(KEYINPUT37), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n748), .B2(new_n424), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n267), .B1(new_n749), .B2(new_n410), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n437), .A2(new_n438), .A3(new_n454), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n517), .A2(new_n267), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n676), .A2(new_n752), .A3(new_n675), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n616), .B(new_n742), .C1(new_n753), .C2(new_n693), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n700), .A2(new_n742), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n661), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n498), .A2(new_n586), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n741), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n505), .A2(G92gat), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n757), .A2(new_n661), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n740), .B2(new_n505), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n740), .A2(new_n766), .A3(new_n505), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n763), .B(new_n765), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G92gat), .B1(new_n740), .B2(new_n505), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n765), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT111), .B1(new_n772), .B2(KEYINPUT52), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n774), .B(new_n763), .C1(new_n771), .C2(new_n765), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n773), .B2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n740), .B2(new_n708), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n503), .A2(new_n583), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n760), .B2(new_n778), .ZN(G1338gat));
  NAND4_X1  g578(.A1(new_n757), .A2(new_n268), .A3(new_n759), .A4(new_n661), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n584), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n782));
  INV_X1    g581(.A(new_n740), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n267), .A2(new_n584), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n781), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n781), .B2(new_n785), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n649), .A2(new_n648), .ZN(new_n791));
  INV_X1    g590(.A(new_n533), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT96), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n530), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n794), .A2(new_n535), .B1(new_n523), .B2(new_n528), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n597), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT10), .B1(new_n796), .B2(KEYINPUT102), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n651), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n650), .ZN(new_n799));
  INV_X1    g598(.A(new_n656), .ZN(new_n800));
  INV_X1    g599(.A(new_n791), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n647), .A4(new_n646), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n800), .A4(new_n803), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n806), .A2(new_n641), .A3(new_n657), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n628), .A2(new_n629), .A3(new_n627), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n620), .B1(new_n619), .B2(new_n622), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n636), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n640), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n661), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n616), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n616), .A2(new_n812), .A3(new_n806), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n807), .A2(new_n657), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n790), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n816), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(new_n616), .A3(new_n812), .A4(new_n806), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n804), .A2(new_n805), .B1(new_n639), .B2(new_n640), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n819), .A2(new_n821), .B1(new_n661), .B2(new_n812), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT114), .B(new_n820), .C1(new_n822), .C2(new_n616), .ZN(new_n823));
  INV_X1    g622(.A(new_n560), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n818), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n560), .A2(new_n642), .A3(new_n617), .A4(new_n660), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n510), .A2(new_n511), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n504), .A2(new_n498), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n641), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n267), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT115), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(new_n503), .A3(new_n829), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n642), .A2(new_n282), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(G1340gat));
  AOI21_X1  g635(.A(G120gat), .B1(new_n830), .B2(new_n661), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n660), .A2(new_n280), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n834), .B2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n274), .A3(new_n560), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n834), .A2(new_n560), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n274), .ZN(G1342gat));
  AOI21_X1  g641(.A(G134gat), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n830), .A2(new_n616), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n834), .A2(new_n616), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n276), .ZN(G1343gat));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n268), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n708), .A2(new_n829), .ZN(new_n850));
  NOR4_X1   g649(.A1(new_n849), .A2(new_n850), .A3(G141gat), .A4(new_n642), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  INV_X1    g651(.A(new_n851), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT58), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n850), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n824), .B1(new_n814), .B2(new_n817), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n826), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .A3(new_n268), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n858), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n268), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(new_n827), .B2(new_n268), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n641), .B(new_n856), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n852), .B(new_n855), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n865), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n865), .B2(G141gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n851), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n849), .A2(new_n850), .ZN(new_n875));
  INV_X1    g674(.A(G148gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n661), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n863), .A2(new_n864), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n850), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n876), .C1(new_n879), .C2(new_n661), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n850), .B(KEYINPUT121), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n827), .A2(KEYINPUT57), .A3(new_n268), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n267), .B1(new_n857), .B2(new_n826), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(new_n661), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n877), .B1(new_n880), .B2(new_n888), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n875), .A2(new_n222), .A3(new_n560), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n878), .A2(new_n824), .A3(new_n850), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n222), .ZN(G1346gat));
  NOR2_X1   g691(.A1(new_n617), .A2(new_n227), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n616), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n879), .A2(new_n893), .B1(new_n894), .B2(new_n227), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n828), .A2(new_n504), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT122), .Z(new_n897));
  AOI21_X1  g696(.A(new_n664), .B1(new_n825), .B2(new_n826), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n641), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n832), .B(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n732), .A2(new_n498), .A3(new_n504), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n642), .A2(new_n353), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  INV_X1    g706(.A(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n833), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G176gat), .B1(new_n909), .B2(new_n660), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n900), .A2(new_n354), .A3(new_n661), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  INV_X1    g711(.A(G183gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n905), .B2(new_n560), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n560), .A2(new_n335), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G183gat), .B1(new_n909), .B2(new_n824), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(new_n916), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n917), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n338), .A3(new_n616), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n833), .A2(new_n616), .A3(new_n908), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(G190gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n924), .B2(G190gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  NAND4_X1  g727(.A1(new_n695), .A2(new_n498), .A3(new_n504), .A4(new_n697), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n886), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n642), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n708), .A2(new_n268), .A3(new_n504), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n898), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n642), .A2(G197gat), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n939), .A2(KEYINPUT124), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT124), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  OR2_X1    g742(.A1(new_n660), .A2(G204gat), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n938), .A2(KEYINPUT62), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n661), .A3(new_n886), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G204gat), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT62), .B1(new_n938), .B2(new_n944), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(G1353gat));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n951), .A3(new_n560), .A4(new_n886), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G211gat), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n929), .A2(new_n930), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n930), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n954), .A2(new_n955), .B1(new_n885), .B2(new_n883), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n951), .B1(new_n956), .B2(new_n560), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n950), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n932), .B2(new_n824), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n952), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n211), .A3(new_n560), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1354gat));
  NOR2_X1   g762(.A1(new_n932), .A2(new_n617), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n616), .A2(new_n212), .ZN(new_n965));
  OAI22_X1  g764(.A1(new_n964), .A2(new_n212), .B1(new_n938), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI221_X1 g767(.A(KEYINPUT127), .B1(new_n938), .B2(new_n965), .C1(new_n964), .C2(new_n212), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1355gat));
endmodule


