//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT88), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT88), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G43gat), .A2(G50gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT15), .B1(new_n212), .B2(new_n207), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n206), .A2(new_n211), .A3(new_n213), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT87), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n217), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n222), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n220), .B1(new_n226), .B2(new_n213), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G22gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G15gat), .ZN(new_n231));
  INV_X1    g030(.A(G15gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT91), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G15gat), .B(G22gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(new_n236), .C1(new_n234), .C2(G1gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G8gat), .ZN(new_n243));
  INV_X1    g042(.A(G8gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT89), .B(new_n220), .C1(new_n226), .C2(new_n213), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n229), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n245), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n239), .B2(new_n241), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT92), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n243), .A2(new_n255), .A3(new_n245), .ZN(new_n256));
  INV_X1    g055(.A(new_n213), .ZN(new_n257));
  NOR4_X1   g056(.A1(KEYINPUT87), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n217), .B2(new_n223), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n221), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT17), .A3(new_n220), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n254), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n248), .B(new_n249), .C1(new_n251), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n249), .B(KEYINPUT13), .Z(new_n266));
  INV_X1    g065(.A(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n246), .B1(new_n229), .B2(new_n247), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT93), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n269), .B(new_n272), .C1(new_n263), .C2(new_n264), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT11), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G197gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT12), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n273), .B(new_n280), .C1(new_n265), .C2(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n290));
  INV_X1    g089(.A(new_n287), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n290), .C1(KEYINPUT26), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT65), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT27), .B(G183gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n297), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(G190gat), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(KEYINPUT65), .A3(new_n294), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n292), .A2(new_n293), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(KEYINPUT64), .A3(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  MUX2_X1   g107(.A(KEYINPUT24), .B(new_n308), .S(new_n293), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n301), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT67), .B(G120gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(G113gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320));
  OR2_X1    g119(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT69), .B1(new_n319), .B2(new_n323), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n316), .A2(G113gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  INV_X1    g129(.A(new_n320), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n326), .A2(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n315), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT72), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n315), .A2(new_n332), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G227gat), .ZN(new_n341));
  INV_X1    g140(.A(G233gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT34), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n333), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT73), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n348));
  INV_X1    g147(.A(new_n346), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n348), .B(new_n349), .C1(new_n337), .C2(new_n333), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n337), .A2(new_n343), .A3(new_n333), .ZN(new_n352));
  XOR2_X1   g151(.A(G15gat), .B(G43gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT70), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT71), .ZN(new_n355));
  XOR2_X1   g154(.A(G71gat), .B(G99gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n352), .B(KEYINPUT32), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n352), .B2(new_n358), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n344), .A2(new_n351), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n359), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n343), .B1(new_n336), .B2(new_n339), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT34), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n365), .A2(new_n366), .B1(new_n347), .B2(new_n350), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n363), .A2(KEYINPUT36), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT36), .B1(new_n363), .B2(new_n368), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT31), .B(G50gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  XOR2_X1   g178(.A(G141gat), .B(G148gat), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT77), .ZN(new_n381));
  XNOR2_X1  g180(.A(G141gat), .B(G148gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT2), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT2), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT78), .B(G155gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(G162gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(new_n386), .ZN(new_n390));
  OAI22_X1  g189(.A1(new_n385), .A2(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G197gat), .B(G204gat), .Z(new_n394));
  INV_X1    g193(.A(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT74), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n396), .B2(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n392), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n391), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n402), .A2(KEYINPUT75), .A3(new_n393), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n393), .B1(new_n402), .B2(KEYINPUT75), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n379), .B1(new_n412), .B2(KEYINPUT82), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT83), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n409), .A3(new_n407), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n391), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n415), .B(new_n416), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n412), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n413), .A2(new_n421), .B1(new_n423), .B2(new_n379), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n378), .B1(new_n424), .B2(G22gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n421), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n379), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n230), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n230), .A3(new_n378), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(G22gat), .A3(new_n375), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n315), .B2(new_n409), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT76), .B1(new_n315), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n435), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n408), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n315), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n436), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n447), .B2(new_n408), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT38), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n442), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n439), .A2(new_n436), .A3(new_n437), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(new_n444), .C1(new_n454), .C2(new_n442), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT85), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(new_n458), .A3(new_n452), .A4(new_n455), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n326), .A2(new_n327), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n330), .A2(new_n331), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(new_n391), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n420), .B2(new_n332), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n420), .A2(new_n332), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n420), .A2(new_n418), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n463), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G57gat), .B(G85gat), .Z(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G1gat), .B(G29gat), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT80), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n481), .B(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n474), .B(new_n477), .C1(new_n471), .C2(new_n468), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n391), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n486), .B2(new_n470), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(new_n473), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n478), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n478), .A2(new_n489), .ZN(new_n491));
  INV_X1    g290(.A(new_n484), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT6), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n494), .B(new_n484), .C1(new_n478), .C2(new_n489), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n490), .A2(new_n493), .B1(new_n495), .B2(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n455), .A2(new_n452), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n446), .A2(new_n436), .A3(new_n408), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n441), .B2(new_n408), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n444), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT38), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n452), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n453), .B(new_n502), .C1(new_n454), .C2(new_n442), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n492), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n460), .A2(new_n496), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n474), .B1(new_n472), .B2(new_n477), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n470), .A3(new_n474), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT39), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n484), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n510), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n511), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(KEYINPUT40), .A3(new_n484), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n491), .A2(new_n492), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n503), .A2(KEYINPUT30), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n499), .B2(new_n502), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n453), .B1(new_n454), .B2(new_n442), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n452), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n516), .A2(new_n519), .A3(new_n520), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n434), .B1(new_n508), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n495), .B1(new_n493), .B2(new_n490), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n433), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n372), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n494), .A3(new_n490), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n505), .ZN(new_n533));
  INV_X1    g332(.A(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n364), .A2(new_n367), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n364), .A2(new_n367), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n433), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT35), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n363), .A2(new_n368), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n426), .A2(G22gat), .A3(new_n427), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n425), .A2(new_n429), .B1(new_n543), .B2(new_n375), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n544), .B2(new_n431), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n491), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n492), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n532), .A2(new_n507), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n525), .ZN(new_n548));
  INV_X1    g347(.A(new_n521), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT35), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n285), .B1(new_n531), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n555), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n243), .B(new_n245), .C1(new_n566), .C2(new_n565), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT94), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n579), .A3(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G134gat), .B(G162gat), .Z(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G99gat), .B(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n592), .B1(new_n589), .B2(new_n591), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n587), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n589), .A2(new_n591), .ZN(new_n602));
  INV_X1    g401(.A(new_n592), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(new_n586), .A3(new_n593), .A4(new_n597), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n601), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n261), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT89), .B1(new_n260), .B2(new_n220), .ZN(new_n609));
  INV_X1    g408(.A(new_n247), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n611), .B2(new_n250), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n600), .A2(new_n605), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT96), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n600), .A2(new_n605), .A3(new_n601), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n229), .A2(new_n614), .A3(new_n247), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n585), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n617), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n611), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n229), .A2(new_n247), .A3(new_n250), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n261), .C1(new_n607), .C2(new_n606), .ZN(new_n626));
  INV_X1    g425(.A(new_n585), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n619), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n621), .B1(new_n619), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n584), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n612), .A2(new_n618), .A3(new_n585), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n627), .B1(new_n624), .B2(new_n626), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n620), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n628), .A3(new_n621), .ZN(new_n635));
  INV_X1    g434(.A(new_n584), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n583), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n600), .A2(new_n565), .A3(new_n605), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n565), .B1(new_n600), .B2(new_n605), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n641), .B2(new_n642), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n565), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n614), .A2(new_n615), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT97), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT98), .B1(new_n661), .B2(new_n644), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n654), .B2(new_n656), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT98), .B(new_n644), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n652), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n657), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n644), .B(KEYINPUT99), .Z(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n650), .B1(new_n671), .B2(new_n646), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n667), .A2(new_n673), .A3(KEYINPUT100), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n644), .B1(new_n663), .B2(new_n664), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n651), .B1(new_n678), .B2(new_n665), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n640), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n553), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n533), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n238), .ZN(G1324gat));
  INV_X1    g484(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n526), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G8gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g490(.A(new_n689), .B(KEYINPUT42), .S(new_n691), .Z(G1325gat));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n369), .B2(new_n370), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT36), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n541), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n363), .A2(KEYINPUT36), .A3(new_n368), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(KEYINPUT101), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G15gat), .B1(new_n683), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n538), .A2(new_n232), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n683), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n683), .A2(new_n433), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NOR3_X1   g504(.A1(new_n583), .A2(new_n639), .A3(new_n681), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n533), .A2(G29gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n553), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT35), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n526), .B1(new_n532), .B2(new_n505), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n545), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n542), .A2(new_n377), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n424), .A2(G22gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n432), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n431), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n550), .B(new_n538), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n532), .A2(new_n507), .A3(new_n546), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT102), .B1(new_n712), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n540), .A2(new_n721), .A3(new_n551), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n457), .A2(new_n501), .A3(new_n503), .A4(new_n459), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n527), .B1(new_n547), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n530), .B1(new_n724), .B2(new_n433), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n720), .B(new_n722), .C1(new_n371), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n726), .B2(new_n638), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n638), .A2(KEYINPUT44), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n531), .B2(new_n552), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n583), .A2(new_n681), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n284), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n727), .A2(new_n533), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n709), .B1(new_n732), .B2(new_n215), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n709), .B(KEYINPUT103), .C1(new_n732), .C2(new_n215), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1328gat));
  NAND2_X1  g536(.A1(new_n553), .A2(new_n706), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n526), .A2(new_n216), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT46), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT104), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n727), .A2(new_n534), .A3(new_n729), .A4(new_n731), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n742), .C1(new_n216), .C2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(G43gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n553), .A2(new_n745), .A3(new_n538), .A4(new_n706), .ZN(new_n746));
  NOR4_X1   g545(.A1(new_n727), .A2(new_n699), .A3(new_n729), .A4(new_n731), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n745), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n727), .A2(new_n372), .A3(new_n729), .A4(new_n731), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n745), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT106), .B(new_n751), .C1(new_n752), .C2(new_n745), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n755), .A3(new_n756), .ZN(G1330gat));
  NOR2_X1   g556(.A1(new_n433), .A2(G50gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n553), .A2(new_n706), .A3(new_n758), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n727), .A2(new_n433), .A3(new_n729), .A4(new_n731), .ZN(new_n760));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT48), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n759), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n720), .A2(new_n722), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n725), .A2(new_n371), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n638), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n729), .ZN(new_n771));
  INV_X1    g570(.A(new_n731), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n770), .A2(new_n434), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n765), .B1(new_n773), .B2(G50gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(KEYINPUT107), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n764), .A2(new_n776), .ZN(G1331gat));
  INV_X1    g576(.A(new_n681), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n640), .A2(new_n284), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n726), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n529), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT109), .B(G57gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  NAND2_X1  g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n526), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n783), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT111), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n782), .A2(new_n792), .A3(new_n783), .A4(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT110), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n794), .B(new_n796), .ZN(G1333gat));
  INV_X1    g596(.A(new_n699), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n782), .A2(G71gat), .A3(new_n798), .A4(new_n783), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n782), .A2(new_n538), .A3(new_n783), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(G71gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n434), .A3(new_n783), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g603(.A1(new_n583), .A2(new_n284), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT112), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n726), .A2(new_n638), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n726), .A2(KEYINPUT51), .A3(new_n638), .A4(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n811), .A2(new_n595), .A3(new_n529), .A4(new_n681), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n806), .A2(new_n681), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n770), .A2(new_n771), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n533), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1336gat));
  NAND2_X1  g615(.A1(new_n526), .A2(new_n596), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n681), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n770), .A2(new_n526), .A3(new_n771), .A4(new_n813), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n822));
  OR2_X1    g621(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n823));
  AND4_X1   g622(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n820), .A2(G92gat), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n819), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(G1337gat));
  INV_X1    g626(.A(G99gat), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n814), .A2(new_n828), .A3(new_n699), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n538), .A3(new_n681), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(G1338gat));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n433), .A2(new_n778), .A3(G106gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G106gat), .B1(new_n814), .B2(new_n433), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n837), .B(new_n834), .C1(new_n835), .C2(new_n832), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1339gat));
  NAND4_X1  g640(.A1(new_n583), .A2(new_n285), .A3(new_n639), .A4(new_n778), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n668), .B2(new_n669), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n678), .B2(new_n665), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n650), .B1(new_n670), .B2(new_n845), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n280), .ZN(new_n852));
  INV_X1    g651(.A(new_n262), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n267), .B1(new_n853), .B2(new_n625), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n267), .A2(new_n268), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n854), .A2(new_n249), .B1(new_n855), .B2(new_n266), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n271), .A2(new_n852), .B1(new_n278), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n638), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n846), .B1(new_n662), .B2(new_n666), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n849), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n667), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT100), .B1(new_n667), .B2(new_n673), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n679), .A2(new_n675), .A3(new_n672), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n284), .A2(new_n860), .A3(new_n851), .A4(new_n667), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(new_n639), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n583), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n638), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT115), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n843), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n533), .A3(new_n539), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n534), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n284), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(G113gat), .ZN(G1340gat));
  NOR2_X1   g677(.A1(new_n875), .A2(new_n778), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n318), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n316), .B2(new_n879), .ZN(G1341gat));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n583), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g682(.A1(new_n639), .A2(new_n526), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(G134gat), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(G134gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n433), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n894), .A3(new_n849), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT116), .B1(new_n848), .B2(new_n850), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT55), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n284), .A2(new_n860), .A3(new_n667), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n865), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n862), .B1(new_n899), .B2(new_n639), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n893), .B1(new_n900), .B2(new_n583), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n842), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n900), .A2(new_n893), .A3(new_n583), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n892), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND4_X1   g703(.A1(new_n284), .A2(new_n860), .A3(new_n851), .A4(new_n667), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n271), .A2(new_n852), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n856), .A2(new_n278), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n674), .B2(new_n680), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n639), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n862), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n869), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n583), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n872), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n842), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n434), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n904), .A2(KEYINPUT118), .B1(new_n916), .B2(new_n891), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n918), .B(new_n892), .C1(new_n902), .C2(new_n903), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n371), .A2(new_n533), .A3(new_n526), .ZN(new_n921));
  INV_X1    g720(.A(G141gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n285), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n699), .A2(new_n434), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT119), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(new_n915), .A3(new_n529), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n534), .A3(new_n284), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n922), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT58), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n924), .A2(KEYINPUT58), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1344gat));
  NOR2_X1   g733(.A1(new_n778), .A2(G148gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n534), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT120), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT57), .B1(new_n873), .B2(new_n433), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n842), .B1(new_n900), .B2(new_n583), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n891), .A3(new_n434), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n681), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n921), .B(KEYINPUT121), .Z(new_n943));
  OR2_X1    g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n938), .B1(new_n944), .B2(G148gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n938), .A2(G148gat), .ZN(new_n946));
  INV_X1    g745(.A(new_n921), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n917), .B2(new_n919), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n681), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n937), .B1(new_n945), .B2(new_n949), .ZN(G1345gat));
  INV_X1    g749(.A(new_n388), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n913), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n920), .A2(new_n921), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n873), .A2(new_n533), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n954), .A2(new_n534), .A3(new_n583), .A4(new_n926), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT122), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n927), .A2(new_n957), .A3(new_n534), .A4(new_n583), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT123), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n953), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1346gat));
  INV_X1    g763(.A(G162gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n927), .A2(new_n965), .A3(new_n884), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT124), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n948), .A2(new_n638), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n965), .ZN(G1347gat));
  NOR2_X1   g768(.A1(new_n529), .A2(new_n534), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n873), .A2(new_n539), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n284), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n681), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g775(.A1(new_n972), .A2(new_n583), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G183gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n978), .B1(new_n297), .B2(new_n977), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n972), .A2(new_n299), .A3(new_n638), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n972), .A2(new_n638), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n983), .B2(G190gat), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT61), .B(new_n299), .C1(new_n972), .C2(new_n638), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g787(.A(KEYINPUT125), .B(new_n981), .C1(new_n984), .C2(new_n985), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1351gat));
  NAND4_X1  g789(.A1(new_n915), .A2(new_n434), .A3(new_n699), .A4(new_n970), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n991), .A2(new_n285), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n798), .A2(new_n971), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n433), .B1(new_n914), .B2(new_n842), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n941), .B(new_n993), .C1(new_n994), .C2(new_n891), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n284), .A2(G197gat), .ZN(new_n996));
  OAI22_X1  g795(.A1(new_n992), .A2(G197gat), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT126), .ZN(G1352gat));
  NOR3_X1   g797(.A1(new_n991), .A2(G204gat), .A3(new_n778), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g799(.A(new_n993), .ZN(new_n1001));
  OAI21_X1  g800(.A(G204gat), .B1(new_n942), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1353gat));
  OR3_X1    g802(.A1(new_n991), .A2(G211gat), .A3(new_n913), .ZN(new_n1004));
  OAI211_X1 g803(.A(KEYINPUT63), .B(G211gat), .C1(new_n995), .C2(new_n913), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n939), .A2(new_n583), .A3(new_n941), .A4(new_n993), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1007), .B2(G211gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1004), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n1011), .B(new_n1004), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1010), .A2(new_n1012), .ZN(G1354gat));
  OAI21_X1  g812(.A(G218gat), .B1(new_n995), .B2(new_n639), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n639), .A2(G218gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1014), .B1(new_n991), .B2(new_n1015), .ZN(G1355gat));
endmodule


