

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795;

  AND2_X1 U368 ( .A1(n645), .A2(n365), .ZN(n393) );
  NAND2_X1 U369 ( .A1(n592), .A2(n591), .ZN(n716) );
  AND2_X1 U370 ( .A1(n665), .A2(n664), .ZN(n347) );
  NOR2_X1 U371 ( .A1(n404), .A2(n402), .ZN(n407) );
  NAND2_X1 U372 ( .A1(n391), .A2(n390), .ZN(n404) );
  XNOR2_X2 U373 ( .A(G137), .B(KEYINPUT5), .ZN(n521) );
  XNOR2_X2 U374 ( .A(n534), .B(n533), .ZN(n779) );
  XNOR2_X2 U375 ( .A(n449), .B(n448), .ZN(n618) );
  XNOR2_X2 U376 ( .A(n616), .B(n419), .ZN(n578) );
  OR2_X1 U377 ( .A1(n354), .A2(n431), .ZN(n430) );
  XNOR2_X1 U378 ( .A(G110), .B(G107), .ZN(n423) );
  XNOR2_X1 U379 ( .A(n620), .B(n619), .ZN(n715) );
  NAND2_X1 U380 ( .A1(n434), .A2(n430), .ZN(n560) );
  XNOR2_X1 U381 ( .A(n509), .B(n508), .ZN(n625) );
  XNOR2_X1 U382 ( .A(n423), .B(G104), .ZN(n772) );
  NAND2_X1 U383 ( .A1(n629), .A2(n628), .ZN(n631) );
  AND2_X1 U384 ( .A1(n409), .A2(n600), .ZN(n602) );
  XNOR2_X1 U385 ( .A(n637), .B(KEYINPUT32), .ZN(n443) );
  AND2_X1 U386 ( .A1(n439), .A2(n438), .ZN(n350) );
  XNOR2_X1 U387 ( .A(n565), .B(n564), .ZN(n702) );
  NAND2_X1 U388 ( .A1(n441), .A2(n442), .ZN(n438) );
  NOR2_X1 U389 ( .A1(n742), .A2(n741), .ZN(n581) );
  NOR2_X1 U390 ( .A1(n589), .A2(n357), .ZN(n449) );
  XNOR2_X1 U391 ( .A(n593), .B(KEYINPUT111), .ZN(n743) );
  NAND2_X1 U392 ( .A1(n585), .A2(n586), .ZN(n713) );
  INV_X1 U393 ( .A(n625), .ZN(n558) );
  AND2_X1 U394 ( .A1(n436), .A2(n435), .ZN(n434) );
  XNOR2_X1 U395 ( .A(n406), .B(n693), .ZN(n695) );
  XNOR2_X1 U396 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U397 ( .A(n547), .B(n546), .ZN(n694) );
  NAND2_X1 U398 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U399 ( .A(n444), .B(n774), .ZN(n547) );
  XNOR2_X1 U400 ( .A(n772), .B(KEYINPUT77), .ZN(n398) );
  XNOR2_X1 U401 ( .A(n782), .B(n490), .ZN(n496) );
  XNOR2_X1 U402 ( .A(n543), .B(n545), .ZN(n445) );
  XNOR2_X1 U403 ( .A(n424), .B(G119), .ZN(n447) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n649) );
  INV_X2 U405 ( .A(G953), .ZN(n785) );
  XNOR2_X1 U406 ( .A(G146), .B(KEYINPUT4), .ZN(n781) );
  NAND2_X1 U407 ( .A1(n385), .A2(n348), .ZN(n349) );
  INV_X1 U408 ( .A(n402), .ZN(n348) );
  NOR2_X1 U409 ( .A1(n349), .A2(n404), .ZN(n368) );
  NOR2_X2 U410 ( .A1(n425), .A2(n358), .ZN(n408) );
  NOR2_X1 U411 ( .A1(n694), .A2(n426), .ZN(n425) );
  NAND2_X1 U412 ( .A1(n439), .A2(n438), .ZN(n747) );
  NAND2_X1 U413 ( .A1(n434), .A2(n430), .ZN(n351) );
  NAND2_X1 U414 ( .A1(n408), .A2(n428), .ZN(n370) );
  NOR2_X1 U415 ( .A1(n352), .A2(n657), .ZN(n376) );
  NAND2_X1 U416 ( .A1(n363), .A2(n608), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n370), .B(n573), .ZN(n353) );
  XNOR2_X2 U418 ( .A(n416), .B(KEYINPUT90), .ZN(n657) );
  XNOR2_X1 U419 ( .A(n370), .B(n573), .ZN(n739) );
  XNOR2_X1 U420 ( .A(n779), .B(n397), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n779), .B(n397), .ZN(n685) );
  NAND2_X1 U422 ( .A1(n625), .A2(n561), .ZN(n722) );
  XNOR2_X2 U423 ( .A(n546), .B(n538), .ZN(n397) );
  INV_X1 U424 ( .A(n415), .ZN(n493) );
  NAND2_X1 U425 ( .A1(n433), .A2(n432), .ZN(n431) );
  INV_X1 U426 ( .A(G146), .ZN(n490) );
  NOR2_X1 U427 ( .A1(n618), .A2(n557), .ZN(n395) );
  XNOR2_X1 U428 ( .A(KEYINPUT73), .B(G137), .ZN(n532) );
  NAND2_X1 U429 ( .A1(KEYINPUT68), .A2(n388), .ZN(n383) );
  NAND2_X1 U430 ( .A1(n364), .A2(KEYINPUT88), .ZN(n384) );
  XNOR2_X1 U431 ( .A(n781), .B(G101), .ZN(n535) );
  XNOR2_X1 U432 ( .A(KEYINPUT24), .B(KEYINPUT87), .ZN(n499) );
  XNOR2_X1 U433 ( .A(G119), .B(KEYINPUT23), .ZN(n500) );
  XOR2_X1 U434 ( .A(KEYINPUT106), .B(KEYINPUT7), .Z(n466) );
  XNOR2_X1 U435 ( .A(G107), .B(KEYINPUT105), .ZN(n465) );
  XOR2_X1 U436 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n468) );
  NAND2_X1 U437 ( .A1(n427), .A2(n649), .ZN(n426) );
  NAND2_X1 U438 ( .A1(n415), .A2(G234), .ZN(n512) );
  INV_X1 U439 ( .A(G134), .ZN(n457) );
  XNOR2_X1 U440 ( .A(G122), .B(G104), .ZN(n484) );
  XNOR2_X1 U441 ( .A(G113), .B(G143), .ZN(n486) );
  XNOR2_X1 U442 ( .A(n482), .B(n412), .ZN(n411) );
  INV_X1 U443 ( .A(G131), .ZN(n412) );
  XNOR2_X1 U444 ( .A(n456), .B(n455), .ZN(n454) );
  INV_X1 U445 ( .A(KEYINPUT28), .ZN(n455) );
  XNOR2_X1 U446 ( .A(n492), .B(n413), .ZN(n591) );
  XNOR2_X1 U447 ( .A(n414), .B(KEYINPUT13), .ZN(n413) );
  INV_X1 U448 ( .A(G475), .ZN(n414) );
  NOR2_X1 U449 ( .A1(n793), .A2(n794), .ZN(n583) );
  XNOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n462) );
  NAND2_X1 U451 ( .A1(n401), .A2(n356), .ZN(n390) );
  AND2_X1 U452 ( .A1(n643), .A2(n356), .ZN(n400) );
  INV_X1 U453 ( .A(KEYINPUT88), .ZN(n388) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n451) );
  NAND2_X1 U455 ( .A1(n364), .A2(n388), .ZN(n387) );
  NAND2_X1 U456 ( .A1(KEYINPUT68), .A2(KEYINPUT88), .ZN(n386) );
  INV_X1 U457 ( .A(n549), .ZN(n427) );
  INV_X1 U458 ( .A(G469), .ZN(n433) );
  NAND2_X1 U459 ( .A1(G902), .A2(G469), .ZN(n435) );
  BUF_X1 U460 ( .A(G237), .Z(n415) );
  XNOR2_X1 U461 ( .A(KEYINPUT79), .B(KEYINPUT100), .ZN(n523) );
  XNOR2_X1 U462 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n545) );
  NAND2_X1 U463 ( .A1(n380), .A2(n377), .ZN(n374) );
  NOR2_X1 U464 ( .A1(n378), .A2(n366), .ZN(n377) );
  INV_X1 U465 ( .A(n363), .ZN(n378) );
  NOR2_X1 U466 ( .A1(n720), .A2(n658), .ZN(n381) );
  INV_X1 U467 ( .A(n722), .ZN(n609) );
  XNOR2_X1 U468 ( .A(n504), .B(n503), .ZN(n662) );
  XNOR2_X1 U469 ( .A(n496), .B(n495), .ZN(n504) );
  XNOR2_X1 U470 ( .A(KEYINPUT107), .B(KEYINPUT9), .ZN(n467) );
  XNOR2_X1 U471 ( .A(G116), .B(G122), .ZN(n471) );
  XNOR2_X1 U472 ( .A(G140), .B(KEYINPUT82), .ZN(n537) );
  NOR2_X1 U473 ( .A1(n519), .A2(n713), .ZN(n596) );
  INV_X1 U474 ( .A(KEYINPUT114), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U476 ( .A(KEYINPUT110), .ZN(n478) );
  INV_X1 U477 ( .A(KEYINPUT0), .ZN(n448) );
  XNOR2_X1 U478 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U479 ( .A(KEYINPUT16), .B(G122), .ZN(n541) );
  XNOR2_X1 U480 ( .A(n411), .B(n483), .ZN(n489) );
  NOR2_X1 U481 ( .A1(n785), .A2(G952), .ZN(n697) );
  NOR2_X1 U482 ( .A1(n588), .A2(n587), .ZN(n710) );
  AND2_X1 U483 ( .A1(n609), .A2(KEYINPUT115), .ZN(n355) );
  OR2_X1 U484 ( .A1(n647), .A2(n646), .ZN(n356) );
  NAND2_X1 U485 ( .A1(n548), .A2(G214), .ZN(n738) );
  NAND2_X1 U486 ( .A1(n556), .A2(n721), .ZN(n357) );
  AND2_X1 U487 ( .A1(n549), .A2(n655), .ZN(n358) );
  AND2_X1 U488 ( .A1(n382), .A2(n381), .ZN(n359) );
  INV_X1 U489 ( .A(G902), .ZN(n432) );
  AND2_X1 U490 ( .A1(n609), .A2(n399), .ZN(n360) );
  NOR2_X1 U491 ( .A1(n396), .A2(n418), .ZN(n361) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT1), .Z(n362) );
  OR2_X1 U493 ( .A1(n656), .A2(KEYINPUT68), .ZN(n363) );
  NAND2_X1 U494 ( .A1(n656), .A2(KEYINPUT68), .ZN(n364) );
  OR2_X1 U495 ( .A1(n653), .A2(n652), .ZN(n365) );
  AND2_X1 U496 ( .A1(n384), .A2(n383), .ZN(n366) );
  NAND2_X1 U497 ( .A1(n649), .A2(n648), .ZN(n367) );
  INV_X1 U498 ( .A(n657), .ZN(n382) );
  XNOR2_X1 U499 ( .A(n553), .B(n552), .ZN(n589) );
  NAND2_X1 U500 ( .A1(n595), .A2(n738), .ZN(n553) );
  AND2_X1 U501 ( .A1(n460), .A2(n458), .ZN(n437) );
  INV_X1 U502 ( .A(n590), .ZN(n453) );
  OR2_X1 U503 ( .A1(n610), .A2(KEYINPUT115), .ZN(n461) );
  AND2_X1 U504 ( .A1(n624), .A2(n623), .ZN(n635) );
  AND2_X1 U505 ( .A1(n458), .A2(n612), .ZN(n442) );
  BUF_X1 U506 ( .A(n711), .Z(n369) );
  NAND2_X1 U507 ( .A1(n453), .A2(n452), .ZN(n711) );
  XNOR2_X1 U508 ( .A(n429), .B(n544), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n444) );
  NAND2_X1 U510 ( .A1(n408), .A2(n428), .ZN(n595) );
  NAND2_X1 U511 ( .A1(n644), .A2(n643), .ZN(n405) );
  NAND2_X1 U512 ( .A1(n572), .A2(n371), .ZN(n575) );
  AND2_X1 U513 ( .A1(n571), .A2(n353), .ZN(n371) );
  INV_X1 U514 ( .A(n589), .ZN(n452) );
  NOR2_X2 U515 ( .A1(G902), .A2(n676), .ZN(n481) );
  NAND2_X1 U516 ( .A1(n403), .A2(n367), .ZN(n402) );
  NOR2_X1 U517 ( .A1(G953), .A2(G237), .ZN(n372) );
  NOR2_X2 U518 ( .A1(G953), .A2(G237), .ZN(n520) );
  NOR2_X2 U519 ( .A1(n657), .A2(n720), .ZN(n654) );
  NAND2_X1 U520 ( .A1(n373), .A2(n379), .ZN(n661) );
  NAND2_X1 U521 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U522 ( .A1(n368), .A2(n376), .ZN(n375) );
  NAND2_X1 U523 ( .A1(n359), .A2(n765), .ZN(n379) );
  NAND2_X1 U524 ( .A1(n654), .A2(n407), .ZN(n380) );
  NAND2_X1 U525 ( .A1(n382), .A2(n608), .ZN(n784) );
  XNOR2_X1 U526 ( .A(n389), .B(n422), .ZN(n421) );
  NAND2_X1 U527 ( .A1(n747), .A2(n613), .ZN(n389) );
  AND2_X1 U528 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U529 ( .A1(n393), .A2(n405), .ZN(n391) );
  NAND2_X1 U530 ( .A1(n640), .A2(n639), .ZN(n644) );
  XNOR2_X1 U531 ( .A(n392), .B(KEYINPUT47), .ZN(n601) );
  NOR2_X2 U532 ( .A1(n711), .A2(n743), .ZN(n392) );
  NAND2_X1 U533 ( .A1(n578), .A2(n577), .ZN(n456) );
  NAND2_X1 U534 ( .A1(n578), .A2(n738), .ZN(n568) );
  XNOR2_X1 U535 ( .A(n394), .B(n451), .ZN(n417) );
  NAND2_X1 U536 ( .A1(n604), .A2(n603), .ZN(n394) );
  XNOR2_X1 U537 ( .A(n395), .B(KEYINPUT22), .ZN(n624) );
  BUF_X1 U538 ( .A(n578), .Z(n396) );
  NAND2_X1 U539 ( .A1(n454), .A2(n579), .ZN(n590) );
  NOR2_X1 U540 ( .A1(n666), .A2(KEYINPUT44), .ZN(n632) );
  XNOR2_X2 U541 ( .A(n398), .B(n535), .ZN(n546) );
  XNOR2_X2 U542 ( .A(n528), .B(G131), .ZN(n534) );
  XNOR2_X2 U543 ( .A(n429), .B(n457), .ZN(n528) );
  NAND2_X1 U544 ( .A1(n610), .A2(n360), .ZN(n617) );
  INV_X1 U545 ( .A(n616), .ZN(n399) );
  XNOR2_X2 U546 ( .A(n560), .B(n362), .ZN(n610) );
  NAND2_X1 U547 ( .A1(n400), .A2(n644), .ZN(n403) );
  INV_X1 U548 ( .A(n645), .ZN(n401) );
  NAND2_X1 U549 ( .A1(n405), .A2(n645), .ZN(n660) );
  XNOR2_X2 U550 ( .A(n631), .B(n630), .ZN(n645) );
  BUF_X1 U551 ( .A(n694), .Z(n406) );
  AND2_X1 U552 ( .A1(n601), .A2(n410), .ZN(n409) );
  INV_X1 U553 ( .A(n710), .ZN(n410) );
  NAND2_X1 U554 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U555 ( .A1(n417), .A2(n606), .ZN(n416) );
  INV_X1 U556 ( .A(n558), .ZN(n418) );
  XNOR2_X2 U557 ( .A(n420), .B(n615), .ZN(n666) );
  NAND2_X1 U558 ( .A1(n421), .A2(n614), .ZN(n420) );
  INV_X1 U559 ( .A(KEYINPUT34), .ZN(n422) );
  XNOR2_X2 U560 ( .A(G116), .B(KEYINPUT76), .ZN(n424) );
  NAND2_X1 U561 ( .A1(n635), .A2(n636), .ZN(n637) );
  NAND2_X1 U562 ( .A1(n694), .A2(n549), .ZN(n428) );
  XNOR2_X2 U563 ( .A(n464), .B(n463), .ZN(n429) );
  NAND2_X1 U564 ( .A1(n685), .A2(G469), .ZN(n436) );
  AND2_X1 U565 ( .A1(n461), .A2(n460), .ZN(n441) );
  NAND2_X1 U566 ( .A1(n437), .A2(n461), .ZN(n440) );
  NAND2_X1 U567 ( .A1(n440), .A2(n611), .ZN(n439) );
  OR2_X2 U568 ( .A1(n667), .A2(G902), .ZN(n531) );
  XNOR2_X2 U569 ( .A(n729), .B(KEYINPUT6), .ZN(n623) );
  NAND2_X1 U570 ( .A1(n443), .A2(n638), .ZN(n642) );
  XNOR2_X1 U571 ( .A(n443), .B(G119), .ZN(G21) );
  XNOR2_X2 U572 ( .A(n542), .B(n541), .ZN(n774) );
  XNOR2_X2 U573 ( .A(n447), .B(n526), .ZN(n542) );
  XNOR2_X2 U574 ( .A(n450), .B(KEYINPUT10), .ZN(n782) );
  XNOR2_X2 U575 ( .A(G125), .B(G140), .ZN(n450) );
  NOR2_X2 U576 ( .A1(n623), .A2(n459), .ZN(n458) );
  NOR2_X1 U577 ( .A1(n609), .A2(KEYINPUT115), .ZN(n459) );
  NAND2_X1 U578 ( .A1(n610), .A2(n355), .ZN(n460) );
  INV_X1 U579 ( .A(n616), .ZN(n729) );
  XNOR2_X2 U580 ( .A(G128), .B(G143), .ZN(n464) );
  XNOR2_X2 U581 ( .A(KEYINPUT66), .B(KEYINPUT85), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n583), .B(n462), .ZN(n604) );
  INV_X1 U583 ( .A(n605), .ZN(n606) );
  INV_X1 U584 ( .A(n532), .ZN(n533) );
  INV_X1 U585 ( .A(G472), .ZN(n530) );
  BUF_X1 U586 ( .A(n667), .Z(n669) );
  INV_X1 U587 ( .A(n697), .ZN(n664) );
  BUF_X1 U588 ( .A(n354), .Z(n687) );
  OR2_X1 U589 ( .A1(n733), .A2(n618), .ZN(n620) );
  XOR2_X1 U590 ( .A(n466), .B(n465), .Z(n470) );
  XNOR2_X1 U591 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U592 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U593 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U594 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n474) );
  NAND2_X1 U595 ( .A1(G234), .A2(n785), .ZN(n473) );
  XNOR2_X1 U596 ( .A(n474), .B(n473), .ZN(n494) );
  NAND2_X1 U597 ( .A1(n494), .A2(G217), .ZN(n475) );
  XNOR2_X1 U598 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U599 ( .A(n528), .B(n477), .ZN(n676) );
  INV_X1 U600 ( .A(G478), .ZN(n479) );
  XNOR2_X2 U601 ( .A(n481), .B(n480), .ZN(n585) );
  XOR2_X1 U602 ( .A(KEYINPUT104), .B(KEYINPUT11), .Z(n483) );
  NAND2_X1 U603 ( .A1(n372), .A2(G214), .ZN(n482) );
  XOR2_X1 U604 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n485) );
  XNOR2_X1 U605 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U606 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U607 ( .A(n489), .B(n488), .ZN(n491) );
  XNOR2_X1 U608 ( .A(n496), .B(n491), .ZN(n680) );
  NOR2_X1 U609 ( .A1(G902), .A2(n680), .ZN(n492) );
  INV_X1 U610 ( .A(n591), .ZN(n586) );
  NAND2_X1 U611 ( .A1(n432), .A2(n493), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n494), .A2(G221), .ZN(n495) );
  XNOR2_X1 U613 ( .A(G110), .B(G128), .ZN(n497) );
  XNOR2_X1 U614 ( .A(n497), .B(KEYINPUT98), .ZN(n498) );
  XNOR2_X1 U615 ( .A(n498), .B(n532), .ZN(n502) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U618 ( .A1(n662), .A2(n432), .ZN(n509) );
  NAND2_X1 U619 ( .A1(n649), .A2(G234), .ZN(n505) );
  XNOR2_X1 U620 ( .A(n505), .B(KEYINPUT20), .ZN(n515) );
  NAND2_X1 U621 ( .A1(n515), .A2(G217), .ZN(n507) );
  XNOR2_X1 U622 ( .A(KEYINPUT81), .B(KEYINPUT25), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U624 ( .A1(G900), .A2(n785), .ZN(n510) );
  NAND2_X1 U625 ( .A1(n510), .A2(G902), .ZN(n511) );
  NAND2_X1 U626 ( .A1(G952), .A2(n785), .ZN(n554) );
  NAND2_X1 U627 ( .A1(n511), .A2(n554), .ZN(n513) );
  XNOR2_X1 U628 ( .A(n512), .B(KEYINPUT14), .ZN(n721) );
  NAND2_X1 U629 ( .A1(n513), .A2(n721), .ZN(n514) );
  XNOR2_X1 U630 ( .A(KEYINPUT86), .B(n514), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G221), .A2(n515), .ZN(n516) );
  XNOR2_X1 U632 ( .A(KEYINPUT21), .B(n516), .ZN(n726) );
  NOR2_X1 U633 ( .A1(n569), .A2(n726), .ZN(n517) );
  NAND2_X1 U634 ( .A1(n558), .A2(n517), .ZN(n518) );
  XNOR2_X1 U635 ( .A(n518), .B(KEYINPUT75), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n738), .A2(n577), .ZN(n519) );
  NAND2_X1 U637 ( .A1(n520), .A2(G210), .ZN(n522) );
  XNOR2_X1 U638 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U639 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U640 ( .A(n525), .B(n535), .ZN(n527) );
  XOR2_X1 U641 ( .A(KEYINPUT3), .B(G113), .Z(n526) );
  XNOR2_X1 U642 ( .A(n527), .B(n542), .ZN(n529) );
  XNOR2_X1 U643 ( .A(n529), .B(n534), .ZN(n667) );
  XNOR2_X2 U644 ( .A(n531), .B(n530), .ZN(n616) );
  INV_X1 U645 ( .A(n623), .ZN(n594) );
  AND2_X1 U646 ( .A1(n596), .A2(n594), .ZN(n539) );
  NAND2_X1 U647 ( .A1(n785), .A2(G227), .ZN(n536) );
  XNOR2_X1 U648 ( .A(n537), .B(n536), .ZN(n538) );
  INV_X1 U649 ( .A(n610), .ZN(n723) );
  NAND2_X1 U650 ( .A1(n539), .A2(n723), .ZN(n540) );
  XOR2_X1 U651 ( .A(KEYINPUT43), .B(n540), .Z(n550) );
  XNOR2_X1 U652 ( .A(G125), .B(KEYINPUT18), .ZN(n544) );
  NAND2_X1 U653 ( .A1(n785), .A2(G224), .ZN(n543) );
  INV_X1 U654 ( .A(n649), .ZN(n655) );
  AND2_X1 U655 ( .A1(n548), .A2(G210), .ZN(n549) );
  NOR2_X1 U656 ( .A1(n550), .A2(n370), .ZN(n605) );
  XOR2_X1 U657 ( .A(G140), .B(n605), .Z(G42) );
  INV_X1 U658 ( .A(KEYINPUT80), .ZN(n551) );
  XNOR2_X1 U659 ( .A(n551), .B(KEYINPUT19), .ZN(n552) );
  XOR2_X1 U660 ( .A(KEYINPUT97), .B(G898), .Z(n767) );
  NOR2_X1 U661 ( .A1(n767), .A2(n785), .ZN(n776) );
  NAND2_X1 U662 ( .A1(n776), .A2(G902), .ZN(n555) );
  NAND2_X1 U663 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U664 ( .A1(n585), .A2(n591), .ZN(n580) );
  XNOR2_X1 U665 ( .A(n726), .B(KEYINPUT99), .ZN(n561) );
  NAND2_X1 U666 ( .A1(n580), .A2(n561), .ZN(n557) );
  AND2_X1 U667 ( .A1(n723), .A2(n361), .ZN(n559) );
  NAND2_X1 U668 ( .A1(n624), .A2(n559), .ZN(n638) );
  XNOR2_X1 U669 ( .A(n638), .B(G110), .ZN(G12) );
  NOR2_X1 U670 ( .A1(n399), .A2(n722), .ZN(n562) );
  NAND2_X1 U671 ( .A1(n351), .A2(n562), .ZN(n563) );
  OR2_X1 U672 ( .A1(n618), .A2(n563), .ZN(n565) );
  INV_X1 U673 ( .A(KEYINPUT101), .ZN(n564) );
  NOR2_X1 U674 ( .A1(n702), .A2(n713), .ZN(n566) );
  XOR2_X1 U675 ( .A(G104), .B(n566), .Z(G6) );
  INV_X1 U676 ( .A(KEYINPUT30), .ZN(n567) );
  XNOR2_X1 U677 ( .A(n568), .B(n567), .ZN(n572) );
  NOR2_X1 U678 ( .A1(n722), .A2(n569), .ZN(n570) );
  AND2_X1 U679 ( .A1(n351), .A2(n570), .ZN(n571) );
  INV_X1 U680 ( .A(KEYINPUT38), .ZN(n573) );
  INV_X1 U681 ( .A(KEYINPUT39), .ZN(n574) );
  XNOR2_X1 U682 ( .A(n575), .B(n574), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n607), .A2(n713), .ZN(n576) );
  XNOR2_X1 U684 ( .A(n576), .B(KEYINPUT40), .ZN(n793) );
  XNOR2_X1 U685 ( .A(n351), .B(KEYINPUT116), .ZN(n579) );
  NAND2_X1 U686 ( .A1(n739), .A2(n738), .ZN(n742) );
  INV_X1 U687 ( .A(n580), .ZN(n741) );
  XNOR2_X1 U688 ( .A(KEYINPUT41), .B(n581), .ZN(n754) );
  NOR2_X1 U689 ( .A1(n590), .A2(n754), .ZN(n582) );
  XNOR2_X1 U690 ( .A(n582), .B(KEYINPUT42), .ZN(n794) );
  INV_X1 U691 ( .A(n584), .ZN(n588) );
  INV_X1 U692 ( .A(n585), .ZN(n592) );
  AND2_X1 U693 ( .A1(n592), .A2(n586), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n614), .A2(n370), .ZN(n587) );
  NAND2_X1 U695 ( .A1(n716), .A2(n713), .ZN(n593) );
  AND2_X1 U696 ( .A1(n370), .A2(n594), .ZN(n597) );
  XNOR2_X1 U697 ( .A(n598), .B(KEYINPUT36), .ZN(n599) );
  XOR2_X1 U698 ( .A(KEYINPUT95), .B(n723), .Z(n633) );
  NOR2_X2 U699 ( .A1(n599), .A2(n633), .ZN(n718) );
  XNOR2_X1 U700 ( .A(n718), .B(KEYINPUT91), .ZN(n600) );
  XNOR2_X1 U701 ( .A(n602), .B(KEYINPUT74), .ZN(n603) );
  OR2_X1 U702 ( .A1(n607), .A2(n716), .ZN(n608) );
  INV_X1 U703 ( .A(n608), .ZN(n720) );
  INV_X1 U704 ( .A(n618), .ZN(n613) );
  XNOR2_X1 U705 ( .A(KEYINPUT78), .B(KEYINPUT33), .ZN(n611) );
  INV_X1 U706 ( .A(n611), .ZN(n612) );
  XNOR2_X1 U707 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n615) );
  NAND2_X1 U708 ( .A1(n666), .A2(KEYINPUT44), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n617), .B(KEYINPUT102), .ZN(n733) );
  INV_X1 U710 ( .A(KEYINPUT31), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n715), .A2(n702), .ZN(n622) );
  INV_X1 U712 ( .A(n743), .ZN(n621) );
  NAND2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n627) );
  XNOR2_X1 U714 ( .A(n418), .B(KEYINPUT112), .ZN(n725) );
  AND2_X1 U715 ( .A1(n723), .A2(n725), .ZN(n626) );
  NAND2_X1 U716 ( .A1(n635), .A2(n626), .ZN(n700) );
  AND2_X1 U717 ( .A1(n627), .A2(n700), .ZN(n628) );
  INV_X1 U718 ( .A(KEYINPUT92), .ZN(n630) );
  XNOR2_X1 U719 ( .A(n632), .B(KEYINPUT71), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n633), .A2(n725), .ZN(n634) );
  XOR2_X1 U721 ( .A(n634), .B(KEYINPUT113), .Z(n636) );
  INV_X1 U722 ( .A(n642), .ZN(n639) );
  INV_X1 U723 ( .A(KEYINPUT44), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  INV_X1 U725 ( .A(KEYINPUT89), .ZN(n648) );
  OR2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U727 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n651) );
  NOR2_X1 U728 ( .A1(n650), .A2(n651), .ZN(n647) );
  INV_X1 U729 ( .A(n651), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n659), .A2(KEYINPUT89), .ZN(n646) );
  NOR2_X1 U731 ( .A1(n650), .A2(n659), .ZN(n653) );
  NOR2_X1 U732 ( .A1(n651), .A2(KEYINPUT89), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n655), .A2(KEYINPUT2), .ZN(n656) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n765) );
  XNOR2_X2 U736 ( .A(n661), .B(KEYINPUT67), .ZN(n691) );
  NAND2_X1 U737 ( .A1(n691), .A2(G217), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n347), .B(KEYINPUT124), .ZN(G66) );
  XOR2_X1 U740 ( .A(n666), .B(G122), .Z(G24) );
  NAND2_X1 U741 ( .A1(n691), .A2(G472), .ZN(n671) );
  XNOR2_X1 U742 ( .A(KEYINPUT94), .B(KEYINPUT62), .ZN(n668) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X2 U744 ( .A1(n672), .A2(n697), .ZN(n674) );
  XOR2_X1 U745 ( .A(KEYINPUT96), .B(KEYINPUT63), .Z(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(G57) );
  BUF_X1 U747 ( .A(n691), .Z(n675) );
  NAND2_X1 U748 ( .A1(n675), .A2(G478), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n678), .A2(n697), .ZN(G63) );
  NAND2_X1 U751 ( .A1(n691), .A2(G475), .ZN(n682) );
  XOR2_X1 U752 ( .A(KEYINPUT70), .B(KEYINPUT59), .Z(n679) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X2 U754 ( .A1(n683), .A2(n697), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n684), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U756 ( .A1(n675), .A2(G469), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U760 ( .A1(n690), .A2(n697), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n691), .A2(G210), .ZN(n696) );
  XNOR2_X1 U762 ( .A(KEYINPUT93), .B(KEYINPUT54), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(KEYINPUT55), .ZN(n693) );
  XNOR2_X1 U764 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X2 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U767 ( .A(G101), .B(n700), .Z(n701) );
  XNOR2_X1 U768 ( .A(n701), .B(KEYINPUT117), .ZN(G3) );
  NOR2_X1 U769 ( .A1(n702), .A2(n716), .ZN(n704) );
  XNOR2_X1 U770 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G107), .B(n705), .ZN(G9) );
  NOR2_X1 U773 ( .A1(n369), .A2(n716), .ZN(n709) );
  XOR2_X1 U774 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n707) );
  XNOR2_X1 U775 ( .A(G128), .B(KEYINPUT29), .ZN(n706) );
  XNOR2_X1 U776 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n709), .B(n708), .ZN(G30) );
  XOR2_X1 U778 ( .A(G143), .B(n710), .Z(G45) );
  NOR2_X1 U779 ( .A1(n369), .A2(n713), .ZN(n712) );
  XOR2_X1 U780 ( .A(G146), .B(n712), .Z(G48) );
  NOR2_X1 U781 ( .A1(n713), .A2(n715), .ZN(n714) );
  XOR2_X1 U782 ( .A(G113), .B(n714), .Z(G15) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U784 ( .A(G116), .B(n717), .Z(G18) );
  XNOR2_X1 U785 ( .A(G125), .B(n718), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U787 ( .A(G134), .B(n720), .Z(G36) );
  NAND2_X1 U788 ( .A1(G952), .A2(n721), .ZN(n753) );
  NAND2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U790 ( .A(n724), .B(KEYINPUT50), .ZN(n732) );
  INV_X1 U791 ( .A(n725), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U793 ( .A(n728), .B(KEYINPUT49), .ZN(n730) );
  NOR2_X1 U794 ( .A1(n730), .A2(n399), .ZN(n731) );
  NAND2_X1 U795 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U797 ( .A(n735), .B(KEYINPUT51), .ZN(n736) );
  XNOR2_X1 U798 ( .A(n736), .B(KEYINPUT120), .ZN(n737) );
  NOR2_X1 U799 ( .A1(n754), .A2(n737), .ZN(n750) );
  NOR2_X1 U800 ( .A1(n353), .A2(n738), .ZN(n740) );
  NOR2_X1 U801 ( .A1(n741), .A2(n740), .ZN(n745) );
  NOR2_X1 U802 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U804 ( .A(KEYINPUT121), .B(n746), .Z(n748) );
  NOR2_X1 U805 ( .A1(n748), .A2(n350), .ZN(n749) );
  NOR2_X1 U806 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U807 ( .A(n751), .B(KEYINPUT52), .ZN(n752) );
  NOR2_X1 U808 ( .A1(n753), .A2(n752), .ZN(n756) );
  NOR2_X1 U809 ( .A1(n754), .A2(n350), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U811 ( .A(KEYINPUT122), .B(n757), .Z(n761) );
  INV_X1 U812 ( .A(n784), .ZN(n758) );
  NAND2_X1 U813 ( .A1(n758), .A2(n765), .ZN(n759) );
  XNOR2_X1 U814 ( .A(n759), .B(KEYINPUT2), .ZN(n760) );
  NOR2_X1 U815 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U816 ( .A1(n785), .A2(n762), .ZN(n763) );
  XNOR2_X1 U817 ( .A(n763), .B(KEYINPUT123), .ZN(n764) );
  XNOR2_X1 U818 ( .A(KEYINPUT53), .B(n764), .ZN(G75) );
  NAND2_X1 U819 ( .A1(n765), .A2(n785), .ZN(n771) );
  NAND2_X1 U820 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U821 ( .A(KEYINPUT61), .B(n766), .ZN(n768) );
  NAND2_X1 U822 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U823 ( .A(n769), .B(KEYINPUT125), .Z(n770) );
  AND2_X1 U824 ( .A1(n771), .A2(n770), .ZN(n778) );
  XOR2_X1 U825 ( .A(n772), .B(G101), .Z(n773) );
  XNOR2_X1 U826 ( .A(n774), .B(n773), .ZN(n775) );
  NOR2_X1 U827 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U828 ( .A(n778), .B(n777), .Z(G69) );
  BUF_X1 U829 ( .A(n779), .Z(n780) );
  XOR2_X1 U830 ( .A(n782), .B(n781), .Z(n783) );
  XNOR2_X1 U831 ( .A(n780), .B(n783), .ZN(n787) );
  XNOR2_X1 U832 ( .A(n784), .B(n787), .ZN(n786) );
  NAND2_X1 U833 ( .A1(n786), .A2(n785), .ZN(n792) );
  XNOR2_X1 U834 ( .A(n787), .B(G227), .ZN(n788) );
  NAND2_X1 U835 ( .A1(n788), .A2(G900), .ZN(n789) );
  XNOR2_X1 U836 ( .A(KEYINPUT126), .B(n789), .ZN(n790) );
  NAND2_X1 U837 ( .A1(G953), .A2(n790), .ZN(n791) );
  NAND2_X1 U838 ( .A1(n792), .A2(n791), .ZN(G72) );
  XOR2_X1 U839 ( .A(n793), .B(G131), .Z(G33) );
  XNOR2_X1 U840 ( .A(G137), .B(KEYINPUT127), .ZN(n795) );
  XNOR2_X1 U841 ( .A(n795), .B(n794), .ZN(G39) );
endmodule

