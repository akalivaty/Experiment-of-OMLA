//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT65), .B(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n208), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n220), .A2(new_n227), .A3(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  OR2_X1    g0054(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(G150), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n230), .B2(new_n201), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n229), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n223), .A2(new_n230), .A3(G1), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n267), .B2(new_n265), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n268), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT73), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n259), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT70), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n286), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G223), .B1(G77), .B2(new_n291), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(G1), .A2(G13), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n295), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(G226), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(G200), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n306), .ZN(new_n308));
  OAI211_X1 g0108(.A(G190), .B(new_n308), .C1(new_n294), .C2(new_n297), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n281), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n255), .B(new_n256), .C1(new_n280), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n310), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n278), .B(KEYINPUT73), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT74), .A4(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n298), .B2(new_n306), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n308), .C1(new_n294), .C2(new_n297), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n276), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n311), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n258), .A2(new_n267), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n275), .B2(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(new_n230), .A3(new_n284), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n324), .A2(KEYINPUT79), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT79), .B1(new_n324), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n284), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT80), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n210), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n209), .B2(G58), .ZN(new_n334));
  INV_X1    g0134(.A(G159), .ZN(new_n335));
  INV_X1    g0135(.A(new_n261), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n334), .A2(new_n230), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n323), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n265), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n324), .A2(new_n325), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n339), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n322), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n305), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n285), .B(new_n346), .C1(G223), .C2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n297), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n303), .B1(new_n304), .B2(new_n241), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n315), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n349), .A2(new_n317), .A3(new_n350), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n345), .A2(KEYINPUT18), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  INV_X1    g0156(.A(new_n322), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT79), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n289), .A2(new_n290), .A3(G20), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(KEYINPUT7), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n324), .A2(KEYINPUT79), .A3(new_n325), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n329), .A2(new_n330), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n329), .A2(new_n330), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n209), .ZN(new_n365));
  INV_X1    g0165(.A(new_n337), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT16), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n342), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n265), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n357), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n354), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n356), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n355), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n351), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n349), .B2(new_n350), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n357), .C1(new_n367), .C2(new_n370), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT17), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n209), .A2(new_n230), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n223), .A2(G1), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(KEYINPUT12), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n267), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(KEYINPUT12), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n269), .A2(G68), .A3(new_n272), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n230), .A2(G33), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n336), .A2(new_n266), .B1(new_n393), .B2(new_n202), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n265), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT11), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  OAI211_X1 g0199(.A(G226), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n400));
  OAI211_X1 g0200(.A(G232), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n402));
  AND3_X1   g0202(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n297), .A2(G238), .A3(new_n301), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n303), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n406), .B2(new_n410), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n399), .B(G169), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n410), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n409), .B1(new_n405), .B2(new_n404), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n407), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n399), .A4(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT76), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n412), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT76), .B1(new_n417), .B2(new_n407), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(G179), .A4(new_n418), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n315), .B1(new_n416), .B2(new_n418), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n399), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n398), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(new_n425), .A3(G190), .A4(new_n418), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(G200), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n430), .A2(new_n431), .A3(new_n397), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G244), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n205), .B2(new_n285), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(G238), .B2(new_n292), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n303), .B1(new_n435), .B2(new_n304), .C1(new_n438), .C2(new_n297), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n257), .A2(new_n336), .B1(new_n230), .B2(new_n202), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n393), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n265), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT72), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n202), .B1(new_n271), .B2(G20), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n269), .A2(new_n446), .B1(new_n202), .B2(new_n267), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n440), .B(new_n449), .C1(new_n375), .C2(new_n439), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n439), .A2(new_n315), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n448), .C1(G179), .C2(new_n439), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n320), .A2(new_n382), .A3(new_n434), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n402), .ZN(new_n455));
  NAND3_X1  g0255(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(KEYINPUT19), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT81), .B(G97), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G87), .A2(G107), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n457), .A2(new_n230), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n230), .B(G68), .C1(new_n289), .C2(new_n290), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G97), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n393), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n265), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n442), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n386), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n271), .A2(G33), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n269), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n468), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n467), .A2(KEYINPUT84), .A3(new_n473), .A4(new_n470), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n300), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G250), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n271), .B2(G45), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n297), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n211), .A2(new_n286), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n435), .A2(G1698), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n487), .C1(new_n289), .C2(new_n290), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n297), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT83), .A3(new_n317), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n300), .A2(new_n480), .B1(new_n297), .B2(new_n483), .ZN(new_n494));
  INV_X1    g0294(.A(new_n489), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G238), .A2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n435), .B2(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n497), .B2(new_n285), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(new_n297), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n499), .B2(G179), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n492), .A2(new_n500), .B1(new_n315), .B2(new_n499), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n494), .B(G190), .C1(new_n498), .C2(new_n297), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  INV_X1    g0303(.A(new_n490), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(G190), .A4(new_n494), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n472), .A2(G87), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n467), .A2(new_n470), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(G200), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n478), .A2(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  NOR2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n480), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(G257), .A3(new_n297), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n517), .B1(new_n524), .B2(new_n405), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT5), .B(G41), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n300), .A2(new_n480), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G169), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n405), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n317), .A3(new_n527), .A4(new_n516), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n336), .A2(new_n202), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n364), .B2(G107), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n462), .A2(new_n464), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n205), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n206), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT82), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT6), .B1(new_n458), .B2(G107), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT82), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n543), .A3(G20), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n339), .B1(new_n533), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n386), .A2(G97), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n472), .B2(G97), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n529), .B(new_n531), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n533), .A2(new_n544), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n265), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n530), .A2(new_n375), .A3(new_n527), .A4(new_n516), .ZN(new_n552));
  INV_X1    g0352(.A(new_n527), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n553), .B(new_n517), .C1(new_n524), .C2(new_n405), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n554), .B2(G200), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n555), .A3(new_n547), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n512), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT86), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n512), .A2(new_n549), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n269), .A2(new_n471), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT25), .B1(new_n267), .B2(new_n205), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n562), .A2(new_n205), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT89), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n489), .A2(G20), .B1(new_n569), .B2(KEYINPUT88), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT87), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n230), .B2(G107), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT88), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(KEYINPUT23), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n230), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n285), .A2(KEYINPUT22), .A3(new_n230), .A4(G87), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT88), .B1(new_n569), .B2(KEYINPUT87), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n230), .B2(G107), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n575), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(new_n570), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n572), .A2(new_n574), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n578), .A4(new_n579), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n568), .B1(new_n589), .B2(new_n265), .ZN(new_n590));
  AOI211_X1 g0390(.A(KEYINPUT89), .B(new_n339), .C1(new_n583), .C2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n567), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  MUX2_X1   g0392(.A(G250), .B(G257), .S(G1698), .Z(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n285), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G33), .A2(G294), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n297), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n515), .A2(G264), .A3(new_n297), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n527), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OR3_X1    g0399(.A1(new_n599), .A2(KEYINPUT90), .A3(new_n315), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT90), .B1(new_n599), .B2(new_n315), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(G179), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n375), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(G200), .B2(new_n599), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n567), .C1(new_n590), .C2(new_n591), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n267), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n562), .B2(new_n610), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n523), .A2(new_n230), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n535), .B2(new_n259), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n264), .A2(new_n229), .B1(G20), .B2(new_n610), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n458), .A2(G33), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT20), .B(new_n616), .C1(new_n619), .C2(new_n614), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G303), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n283), .A2(new_n622), .A3(new_n284), .ZN(new_n623));
  MUX2_X1   g0423(.A(G257), .B(G264), .S(G1698), .Z(new_n624));
  OAI211_X1 g0424(.A(new_n405), .B(new_n623), .C1(new_n624), .C2(new_n291), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n515), .A2(G270), .A3(new_n297), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n527), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n609), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n618), .A2(new_n620), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n472), .A2(G116), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n611), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .A4(new_n627), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n625), .A2(new_n527), .A3(new_n626), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G190), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n621), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n632), .A2(G179), .A3(new_n634), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n629), .A2(new_n633), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n454), .A2(new_n561), .A3(new_n608), .A4(new_n639), .ZN(G372));
  OR2_X1    g0440(.A1(new_n452), .A2(new_n432), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n429), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(KEYINPUT95), .A3(new_n429), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n644), .A2(new_n381), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n355), .A2(new_n373), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n311), .B(new_n314), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n319), .ZN(new_n649));
  INV_X1    g0449(.A(new_n454), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n499), .A2(G179), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n315), .B2(new_n499), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n499), .A2(KEYINPUT91), .A3(G200), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT91), .B1(new_n499), .B2(G200), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n478), .A2(new_n652), .B1(new_n510), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n607), .A3(new_n549), .A4(new_n556), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n629), .A2(new_n633), .A3(new_n638), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n589), .A2(new_n265), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n589), .A2(new_n568), .A3(new_n265), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n566), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n603), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT93), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n661), .B1(new_n592), .B2(new_n603), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT93), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n660), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n549), .A2(new_n556), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT92), .A3(new_n607), .A4(new_n657), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n463), .A2(G97), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n260), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT19), .ZN(new_n679));
  AOI21_X1  g0479(.A(G20), .B1(new_n283), .B2(new_n284), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n678), .A2(new_n679), .B1(new_n680), .B2(G68), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n458), .A2(new_n459), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n403), .A2(new_n402), .A3(new_n679), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(G20), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n469), .B1(new_n685), .B2(new_n265), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT84), .B1(new_n686), .B2(new_n473), .ZN(new_n687));
  INV_X1    g0487(.A(new_n477), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n501), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n510), .A2(new_n511), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT26), .B1(new_n691), .B2(new_n549), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n478), .A2(new_n652), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n531), .B1(new_n554), .B2(G169), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n551), .B2(new_n547), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n657), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n551), .A2(new_n547), .ZN(new_n702));
  INV_X1    g0502(.A(new_n694), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n689), .A3(new_n703), .A4(new_n690), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT94), .A3(new_n697), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n673), .A2(new_n675), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n649), .B1(new_n650), .B2(new_n707), .ZN(G369));
  NAND2_X1  g0508(.A1(new_n604), .A2(new_n607), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n384), .A2(new_n230), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(G213), .ZN(new_n713));
  INV_X1    g0513(.A(G343), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n666), .A2(new_n716), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n709), .A2(new_n717), .B1(new_n604), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n632), .A2(new_n715), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n639), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n662), .B2(new_n719), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(G330), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n662), .A2(new_n715), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n608), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n592), .A2(new_n603), .A3(new_n716), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n723), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n225), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n682), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n233), .B2(new_n731), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n604), .A2(new_n607), .A3(new_n639), .A4(new_n716), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n561), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT97), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n599), .A2(new_n634), .A3(G179), .A4(new_n491), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n530), .A2(new_n516), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n739), .B(new_n744), .C1(new_n740), .C2(new_n741), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n599), .A2(new_n491), .A3(G179), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n746), .B(new_n627), .C1(new_n553), .C2(new_n741), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n748), .A2(new_n749), .A3(new_n715), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n748), .B2(new_n715), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n700), .A2(new_n706), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n675), .A2(new_n660), .A3(new_n669), .A4(new_n672), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n757), .B(new_n715), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n698), .A2(new_n699), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT94), .B1(new_n705), .B2(new_n697), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT98), .B1(new_n763), .B2(new_n716), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n756), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n607), .A2(new_n549), .A3(new_n556), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT99), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n766), .A2(new_n668), .A3(new_n767), .A4(new_n657), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT99), .B1(new_n658), .B2(new_n670), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n693), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n696), .B1(new_n657), .B2(new_n695), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n715), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT29), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n755), .B1(new_n765), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n735), .B1(new_n776), .B2(G1), .ZN(G364));
  AOI21_X1  g0577(.A(new_n229), .B1(G20), .B2(new_n315), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n230), .A2(G179), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n285), .B1(new_n782), .B2(G329), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n230), .A2(new_n317), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n784), .B(KEYINPUT101), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n375), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n793), .B2(G322), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n790), .A2(new_n780), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n779), .A2(new_n375), .A3(G200), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n622), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n230), .B1(new_n791), .B2(new_n317), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n785), .A2(new_n375), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(G326), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n797), .A2(new_n801), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n809));
  INV_X1    g0609(.A(new_n805), .ZN(new_n810));
  INV_X1    g0610(.A(G58), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n285), .B1(new_n266), .B2(new_n810), .C1(new_n792), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n796), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G77), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n781), .A2(new_n335), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT32), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(KEYINPUT32), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n787), .A2(new_n340), .B1(new_n204), .B2(new_n802), .ZN(new_n819));
  INV_X1    g0619(.A(G87), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n820), .A2(new_n800), .B1(new_n799), .B2(new_n205), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT103), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n807), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n778), .B1(new_n809), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n223), .A2(G20), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n271), .B1(new_n828), .B2(G45), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n730), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n225), .A2(G355), .A3(new_n285), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n249), .A2(new_n479), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n729), .A2(new_n285), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(G45), .B2(new_n233), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n833), .B1(G116), .B2(new_n225), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(G13), .A2(G33), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(G20), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n778), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n832), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n826), .B1(new_n827), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n827), .B2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n840), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n721), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n721), .A2(G330), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n721), .A2(G330), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n832), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(G396));
  NOR2_X1   g0650(.A1(new_n452), .A2(new_n715), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n450), .B1(new_n449), .B2(new_n716), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n452), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n760), .B2(new_n764), .ZN(new_n855));
  INV_X1    g0655(.A(new_n453), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n763), .A2(new_n856), .A3(new_n716), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n831), .B1(new_n858), .B2(new_n754), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n754), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n778), .A2(new_n838), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT104), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n831), .B1(new_n862), .B2(G77), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G137), .A2(new_n805), .B1(new_n786), .B2(G150), .ZN(new_n864));
  INV_X1    g0664(.A(G143), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n864), .B1(new_n796), .B2(new_n335), .C1(new_n865), .C2(new_n792), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT34), .Z(new_n867));
  OAI22_X1  g0667(.A1(new_n266), .A2(new_n800), .B1(new_n799), .B2(new_n340), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT106), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  INV_X1    g0671(.A(new_n802), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G58), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n291), .B1(new_n782), .B2(G132), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n792), .A2(new_n803), .B1(new_n204), .B2(new_n802), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT105), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n291), .B1(new_n781), .B2(new_n795), .C1(new_n810), .C2(new_n622), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n813), .B2(G116), .ZN(new_n879));
  INV_X1    g0679(.A(new_n800), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n786), .A2(G283), .B1(new_n880), .B2(G107), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(new_n820), .C2(new_n799), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n867), .A2(new_n875), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n863), .B1(new_n883), .B2(new_n778), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n853), .B2(new_n839), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n860), .A2(new_n885), .ZN(G384));
  AOI211_X1 g0686(.A(new_n202), .B(new_n233), .C1(new_n209), .C2(G58), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n340), .A2(G50), .ZN(new_n888));
  OAI211_X1 g0688(.A(G1), .B(new_n223), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT108), .Z(new_n890));
  NAND2_X1  g0690(.A1(new_n540), .A2(new_n543), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  OAI211_X1 g0692(.A(G116), .B(new_n231), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(KEYINPUT36), .ZN(new_n897));
  INV_X1    g0697(.A(new_n775), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n650), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n765), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n900), .A2(new_n649), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT110), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n380), .B1(new_n345), .B2(new_n354), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n713), .B(KEYINPUT109), .Z(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n345), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT37), .B1(new_n371), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n371), .A2(new_n372), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(KEYINPUT110), .A3(new_n910), .A4(new_n380), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n357), .B1(new_n370), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n713), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n372), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n904), .B1(new_n916), .B2(new_n380), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n914), .A2(new_n915), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n382), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n917), .B1(new_n908), .B2(new_n911), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n374), .B2(new_n381), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n398), .A2(new_n715), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n429), .A2(new_n433), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n419), .A2(G169), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT14), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(new_n426), .A3(new_n414), .A4(new_n421), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n398), .B(new_n715), .C1(new_n933), .C2(new_n432), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n453), .B(new_n715), .C1(new_n758), .C2(new_n759), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n928), .B(new_n935), .C1(new_n936), .C2(new_n851), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n647), .A2(new_n906), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n371), .A2(new_n905), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n910), .A2(new_n939), .A3(new_n380), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n908), .A2(new_n911), .B1(KEYINPUT37), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n374), .B2(new_n381), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n924), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n923), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n429), .A2(new_n715), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n923), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n937), .A2(new_n938), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n901), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n736), .B1(new_n558), .B2(new_n560), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n750), .A2(new_n751), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n853), .B(new_n935), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n955), .A3(KEYINPUT40), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n927), .B2(new_n923), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(KEYINPUT40), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n454), .A2(new_n753), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(G330), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n951), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n271), .B2(new_n828), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n951), .A2(new_n962), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n897), .B1(KEYINPUT36), .B2(new_n896), .C1(new_n964), .C2(new_n965), .ZN(G367));
  INV_X1    g0766(.A(new_n776), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n725), .B1(new_n718), .B2(new_n724), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(new_n848), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n757), .B1(new_n707), .B2(new_n715), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n763), .A2(KEYINPUT98), .A3(new_n716), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT29), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n754), .B(new_n969), .C1(new_n972), .C2(new_n898), .ZN(new_n973));
  INV_X1    g0773(.A(new_n723), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n702), .A2(new_n715), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n674), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n695), .A2(new_n715), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n727), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n727), .A2(new_n978), .A3(KEYINPUT44), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n727), .B2(new_n978), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n976), .A2(new_n977), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n985), .A2(new_n725), .A3(KEYINPUT45), .A4(new_n726), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n981), .A2(new_n982), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n974), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT112), .B1(new_n973), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n723), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT112), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n776), .A2(new_n990), .A3(new_n991), .A4(new_n969), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n967), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n730), .B(new_n994), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n829), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n985), .A2(new_n608), .A3(new_n724), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n549), .B1(new_n976), .B2(new_n604), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n998), .A2(KEYINPUT42), .B1(new_n716), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT42), .B2(new_n998), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n509), .A2(new_n715), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n693), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n657), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1001), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n974), .A2(new_n978), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n997), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n835), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n239), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n841), .B1(new_n225), .B2(new_n442), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n831), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n802), .A2(new_n340), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n787), .A2(new_n335), .B1(new_n810), .B2(new_n865), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n799), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(G77), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(G137), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n285), .B1(new_n781), .B2(new_n1020), .C1(new_n811), .C2(new_n800), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n813), .B2(G50), .ZN(new_n1022));
  INV_X1    g0822(.A(G150), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1022), .C1(new_n1023), .C2(new_n792), .ZN(new_n1024));
  INV_X1    g0824(.A(G317), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n291), .B1(new_n781), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G294), .B2(new_n786), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n796), .B2(new_n798), .C1(new_n622), .C2(new_n792), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n880), .A2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT46), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n872), .A2(G107), .B1(new_n1018), .B2(new_n535), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n795), .C2(new_n810), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1034), .B2(new_n778), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1005), .A2(new_n840), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1011), .A2(new_n1037), .ZN(G387));
  OR2_X1    g0838(.A1(new_n718), .A2(new_n845), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n244), .A2(new_n479), .A3(new_n285), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT50), .B1(new_n257), .B2(G50), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n479), .C1(new_n340), .C2(new_n202), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n257), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n291), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n732), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n729), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n841), .B1(new_n205), .B2(new_n225), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n831), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n285), .B1(new_n781), .B2(new_n1023), .C1(new_n202), .C2(new_n800), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n813), .B2(G68), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n805), .A2(G159), .B1(new_n1018), .B2(G97), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n786), .A2(new_n258), .B1(new_n872), .B2(new_n468), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n793), .A2(G50), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n285), .B1(new_n782), .B2(G326), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n802), .A2(new_n798), .B1(new_n800), .B2(new_n803), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G311), .A2(new_n786), .B1(new_n805), .B2(G322), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n796), .B2(new_n622), .C1(new_n1025), .C2(new_n792), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1055), .B1(new_n610), .B2(new_n799), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n778), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n969), .A2(new_n830), .B1(new_n1039), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n973), .A2(new_n730), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n776), .A2(new_n969), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n990), .A2(new_n830), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n253), .A2(new_n1012), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n841), .B1(new_n225), .B2(new_n458), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n831), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n792), .A2(new_n335), .B1(new_n1023), .B2(new_n810), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n802), .A2(new_n202), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n210), .A2(new_n800), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G50), .C2(new_n786), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n285), .B1(new_n781), .B2(new_n865), .C1(new_n820), .C2(new_n799), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n813), .B2(new_n258), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n792), .A2(new_n795), .B1(new_n1025), .B2(new_n810), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  AOI21_X1  g0884(.A(new_n285), .B1(new_n782), .B2(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n205), .B2(new_n799), .C1(new_n796), .C2(new_n803), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n800), .A2(new_n798), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n787), .A2(new_n622), .B1(new_n610), .B2(new_n802), .ZN(new_n1088));
  OR3_X1    g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1082), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1074), .B1(new_n1090), .B2(new_n778), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n985), .B2(new_n845), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1071), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n989), .A2(new_n992), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n731), .B1(new_n973), .B2(new_n988), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(G390));
  NAND4_X1  g0897(.A1(new_n753), .A2(G330), .A3(new_n853), .A4(new_n935), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n923), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT39), .B1(new_n923), .B2(new_n943), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n935), .B1(new_n936), .B2(new_n851), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n947), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n944), .A2(new_n1104), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n770), .A2(new_n773), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n852), .A2(new_n452), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n716), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n851), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1106), .B1(new_n935), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1099), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n935), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n857), .B2(new_n1110), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1115), .A2(new_n947), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n935), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1104), .A3(new_n944), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1118), .A3(new_n1098), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n853), .C1(new_n952), .C2(new_n953), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1114), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1098), .A2(new_n1122), .A3(new_n1110), .A4(new_n1109), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1121), .B(new_n935), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n715), .B1(new_n758), .B2(new_n759), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n851), .B1(new_n1125), .B2(new_n856), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n755), .A2(new_n454), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n900), .A2(new_n1127), .A3(new_n649), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n731), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT116), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1113), .A2(new_n830), .A3(new_n1119), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT113), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1113), .A2(KEYINPUT113), .A3(new_n830), .A4(new_n1119), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n831), .B1(new_n862), .B2(new_n258), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n810), .A2(new_n798), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1077), .B(new_n1139), .C1(G107), .C2(new_n786), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n799), .A2(new_n340), .B1(new_n781), .B2(new_n803), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n813), .B2(new_n535), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n610), .C2(new_n792), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n291), .B1(new_n800), .B2(new_n820), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT115), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n291), .B1(new_n782), .B2(G125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n266), .B2(new_n799), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT114), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n787), .A2(new_n1020), .B1(new_n335), .B2(new_n802), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G128), .B2(new_n805), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n793), .A2(G132), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  NAND2_X1  g0952(.A1(new_n813), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n800), .A2(new_n1023), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1143), .A2(new_n1145), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1138), .B1(new_n1157), .B2(new_n778), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1102), .B2(new_n839), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1132), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(KEYINPUT116), .B(new_n1161), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1131), .B1(new_n1160), .B2(new_n1162), .ZN(G378));
  INV_X1    g0963(.A(KEYINPUT119), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  OAI21_X1  g0965(.A(G330), .B1(new_n957), .B2(KEYINPUT40), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n956), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n276), .A2(new_n915), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n320), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n311), .A2(new_n314), .A3(new_n319), .A4(new_n1168), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1166), .A2(new_n1167), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1176), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n928), .A2(new_n955), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT40), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1185), .B2(new_n956), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n950), .B1(new_n1178), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1177), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n937), .A2(new_n938), .A3(new_n949), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n956), .A3(new_n1181), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1165), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1165), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1116), .A2(new_n1118), .A3(new_n1098), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1098), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n1129), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n900), .A2(new_n649), .A3(new_n1128), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1164), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n731), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1189), .B1(new_n1190), .B2(new_n1188), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT118), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1193), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1127), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n901), .B(new_n1128), .C1(new_n1120), .C2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n1211), .A3(KEYINPUT119), .A4(KEYINPUT57), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1201), .A2(new_n1205), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n799), .A2(new_n811), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n787), .A2(new_n204), .B1(new_n800), .B2(new_n202), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G116), .C2(new_n805), .ZN(new_n1216));
  INV_X1    g1016(.A(G41), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n291), .C1(new_n781), .C2(new_n798), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1016), .B(new_n1218), .C1(new_n793), .C2(G107), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(new_n442), .C2(new_n796), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n291), .A2(new_n1217), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G50), .B1(new_n259), .B2(new_n1217), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1220), .A2(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n793), .B1(new_n813), .B2(G137), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n805), .A2(G125), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n786), .A2(G132), .B1(new_n872), .B2(G150), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n880), .A2(new_n1152), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT117), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1018), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1224), .B1(new_n1221), .B2(new_n1220), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n778), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n832), .B1(new_n266), .B2(new_n861), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n1177), .C2(new_n839), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1202), .B2(new_n830), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1213), .A2(new_n1243), .ZN(G375));
  NAND2_X1  g1044(.A1(new_n1199), .A2(new_n1210), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n995), .A3(new_n1129), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1114), .A2(new_n838), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n831), .B1(new_n862), .B2(G68), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n291), .B(new_n1214), .C1(G128), .C2(new_n782), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n872), .A2(G50), .B1(new_n880), .B2(G159), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G132), .A2(new_n805), .B1(new_n786), .B2(new_n1152), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n792), .B2(new_n1020), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1251), .B1(new_n1252), .B2(new_n1254), .C1(new_n1023), .C2(new_n796), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1252), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n291), .B1(new_n799), .B2(new_n202), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT120), .Z(new_n1258));
  OAI22_X1  g1058(.A1(new_n787), .A2(new_n610), .B1(new_n810), .B2(new_n803), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G97), .B2(new_n880), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n793), .A2(G283), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n813), .A2(G107), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n872), .A2(new_n468), .B1(new_n782), .B2(G303), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1255), .A2(new_n1256), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1248), .B1(new_n1265), .B2(new_n778), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1127), .A2(new_n830), .B1(new_n1247), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1246), .A2(new_n1267), .ZN(G381));
  OR2_X1    g1068(.A1(G393), .A2(G396), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(G384), .A3(G381), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(new_n1011), .A3(new_n1037), .A4(new_n1096), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(KEYINPUT122), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1131), .A2(new_n1137), .A3(new_n1159), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G375), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(KEYINPUT122), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .ZN(G407));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1275), .B2(new_n714), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G407), .A2(new_n1279), .ZN(G409));
  NAND3_X1  g1080(.A1(G378), .A2(new_n1213), .A3(new_n1243), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1242), .B1(new_n1209), .B2(new_n830), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n996), .B2(new_n1203), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1278), .A2(G343), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n1245), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n730), .B1(new_n1289), .B2(new_n1245), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1267), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1267), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1286), .A2(new_n1288), .A3(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1287), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1296), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1306), .A2(new_n1307), .B1(KEYINPUT123), .B2(new_n1297), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1287), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1299), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1297), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1300), .A2(new_n1309), .A3(new_n1310), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G387), .A2(new_n1096), .ZN(new_n1316));
  XOR2_X1   g1116(.A(G393), .B(G396), .Z(new_n1317));
  NAND3_X1  g1117(.A1(new_n1011), .A2(new_n1037), .A3(G390), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1317), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1011), .B2(new_n1037), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1037), .ZN(new_n1322));
  AOI211_X1 g1122(.A(new_n1322), .B(new_n1096), .C1(new_n997), .C2(new_n1010), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1320), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1319), .A2(new_n1324), .A3(KEYINPUT126), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT126), .B1(new_n1319), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1315), .A2(new_n1327), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1304), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1331));
  AOI211_X1 g1131(.A(KEYINPUT123), .B(new_n1305), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1329), .B(new_n1310), .C1(new_n1311), .C2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1298), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT124), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1298), .B2(new_n1336), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1311), .A2(KEYINPUT124), .A3(KEYINPUT63), .A4(new_n1297), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1335), .A2(new_n1337), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1328), .A2(new_n1341), .ZN(G405));
  NAND2_X1  g1142(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT126), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  AND3_X1   g1145(.A1(G378), .A2(new_n1213), .A3(new_n1243), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1274), .B1(new_n1213), .B2(new_n1243), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1297), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1319), .A2(new_n1324), .A3(KEYINPUT126), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1284), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1281), .A3(new_n1296), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1345), .A2(new_n1348), .A3(new_n1349), .A4(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1346), .A2(new_n1347), .A3(new_n1297), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1296), .B1(new_n1350), .B2(new_n1281), .ZN(new_n1356));
  OAI22_X1  g1156(.A1(new_n1355), .A2(new_n1356), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1357), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1354), .A2(new_n1358), .ZN(G402));
endmodule


