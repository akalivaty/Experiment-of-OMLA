//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(new_n456), .B(KEYINPUT68), .Z(G261));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .A3(G137), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  INV_X1    g057(.A(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n478), .A2(new_n475), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(G136), .B2(new_n491), .ZN(G162));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n475), .B1(KEYINPUT70), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n495), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n498), .B2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(new_n493), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n475), .A3(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n467), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(G138), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n512), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n478), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(G138), .B(new_n475), .C1(new_n465), .C2(new_n466), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT4), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n501), .A2(new_n507), .B1(new_n515), .B2(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n526), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT75), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  AND2_X1   g110(.A1(new_n528), .A2(G89), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n523), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(G51), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n520), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(KEYINPUT6), .A2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(KEYINPUT6), .A2(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(KEYINPUT73), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n538), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n535), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n525), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT76), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n523), .A2(new_n528), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n549), .A2(KEYINPUT76), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n553), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  INV_X1    g132(.A(new_n545), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G43), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n525), .ZN(new_n561));
  INV_X1    g136(.A(new_n552), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G81), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g146(.A1(new_n528), .A2(new_n540), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n572), .A2(G53), .A3(G543), .A4(new_n544), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n541), .A2(new_n575), .A3(G53), .A4(new_n544), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n562), .A2(G91), .ZN(new_n578));
  INV_X1    g153(.A(new_n522), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT5), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G65), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n578), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n577), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  INV_X1    g165(.A(G168), .ZN(G286));
  AND3_X1   g166(.A1(new_n541), .A2(G49), .A3(new_n544), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n552), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G288));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n521), .B2(new_n522), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n523), .A2(new_n528), .A3(G86), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n528), .A2(G48), .A3(G543), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n558), .A2(G47), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n525), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n562), .A2(G85), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n552), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n558), .A2(G54), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n525), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n619), .C1(new_n613), .C2(new_n614), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT79), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G321));
  XNOR2_X1  g199(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n589), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G868), .B2(new_n589), .ZN(G280));
  INV_X1    g203(.A(new_n623), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G860), .B2(new_n623), .ZN(G148));
  OAI21_X1  g206(.A(G868), .B1(new_n629), .B2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n478), .A2(new_n472), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n485), .A2(G123), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n642), .C1(new_n643), .C2(new_n490), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT82), .B(G2096), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n639), .A2(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  INV_X1    g244(.A(new_n666), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n664), .B2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(KEYINPUT85), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n664), .B(KEYINPUT17), .Z(new_n674));
  INV_X1    g249(.A(new_n665), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n672), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n666), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n669), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n685));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n682), .A2(new_n683), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n687), .B2(new_n684), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(KEYINPUT87), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT88), .Z(new_n696));
  XOR2_X1   g271(.A(G1981), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n696), .B(new_n701), .Z(G229));
  NOR2_X1   g277(.A1(G16), .A2(G23), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n592), .A2(new_n595), .A3(KEYINPUT91), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT91), .B1(new_n592), .B2(new_n595), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G6), .B(G305), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT90), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n712), .A2(new_n713), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n710), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n715), .A2(G24), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n715), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n485), .A2(G119), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n475), .A2(G107), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n730), .B2(new_n731), .C1(new_n732), .C2(new_n490), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G25), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT89), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT92), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n724), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n722), .A2(new_n723), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT36), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n747), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n565), .B2(G16), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1341), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n759), .B(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G11), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(G11), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n735), .B1(new_n767), .B2(G28), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n765), .B(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n644), .A2(new_n735), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(KEYINPUT97), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n763), .B(new_n772), .C1(KEYINPUT97), .C2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT24), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(KEYINPUT94), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(KEYINPUT94), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n481), .B2(new_n735), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n757), .B(new_n773), .C1(new_n774), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n756), .A2(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n735), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n491), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G128), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n784), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n782), .B(new_n791), .C1(new_n774), .C2(new_n780), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT96), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT95), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT26), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n485), .A2(G129), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n472), .A2(G105), .ZN(new_n799));
  INV_X1    g374(.A(G141), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n490), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n796), .B2(KEYINPUT26), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G32), .B(new_n803), .S(G29), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT27), .B(G1996), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n781), .A2(new_n793), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n715), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n623), .B2(new_n715), .ZN(new_n809));
  INV_X1    g384(.A(G1348), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n715), .A2(G20), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n589), .B2(new_n715), .ZN(new_n814));
  INV_X1    g389(.A(G1956), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G171), .A2(new_n715), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G5), .B2(new_n715), .ZN(new_n819));
  INV_X1    g394(.A(G1961), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n735), .A2(G33), .ZN(new_n822));
  NAND2_X1  g397(.A1(G115), .A2(G2104), .ZN(new_n823));
  INV_X1    g398(.A(G127), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n467), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n475), .B1(new_n825), .B2(KEYINPUT93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT93), .B2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n828));
  NAND2_X1  g403(.A1(G103), .A2(G2104), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(G2105), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n475), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n491), .A2(G139), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n822), .B1(new_n834), .B2(new_n735), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G2072), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n715), .A2(G21), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G168), .B2(new_n715), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n821), .B(new_n836), .C1(G1966), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n735), .A2(G27), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G164), .B2(new_n735), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n838), .A2(G1966), .B1(G2078), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n842), .B1(G2078), .B2(new_n841), .C1(new_n819), .C2(new_n820), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n807), .A2(new_n817), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n754), .A2(new_n844), .ZN(G150));
  INV_X1    g420(.A(G150), .ZN(G311));
  NAND2_X1  g421(.A1(new_n623), .A2(G559), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT38), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n523), .A2(G67), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n525), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n552), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT100), .B(G55), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n851), .A2(KEYINPUT99), .B1(new_n545), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n565), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n848), .B(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n860), .A2(new_n861), .A3(G860), .ZN(new_n862));
  OAI21_X1  g437(.A(G860), .B1(new_n854), .B2(new_n856), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT101), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  OR2_X1    g440(.A1(new_n862), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n733), .B(new_n637), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n485), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n870));
  INV_X1    g445(.A(G142), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n870), .C1(new_n871), .C2(new_n490), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT102), .Z(new_n874));
  INV_X1    g449(.A(new_n789), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n797), .A2(new_n875), .A3(new_n802), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n797), .B2(new_n802), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n505), .A2(new_n493), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n515), .B2(new_n517), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n833), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n834), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(G162), .B(new_n644), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n481), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n884), .A2(new_n885), .A3(new_n873), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(G37), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n874), .A2(new_n885), .A3(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n896), .B(new_n898), .ZN(G395));
  XNOR2_X1  g474(.A(new_n630), .B(new_n858), .ZN(new_n900));
  AND2_X1   g475(.A1(G299), .A2(new_n621), .ZN(new_n901));
  NOR2_X1   g476(.A1(G299), .A2(new_n621), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(KEYINPUT105), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n901), .B2(new_n902), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n900), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n707), .A2(new_n726), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n706), .A2(G290), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT106), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(G305), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(KEYINPUT42), .Z(new_n925));
  AND2_X1   g500(.A1(new_n913), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n913), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G868), .B2(new_n857), .ZN(G295));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n857), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n858), .A2(G168), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n857), .B(new_n564), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G286), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n937), .A3(G171), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G171), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n903), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G301), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(new_n938), .A3(new_n904), .A4(new_n905), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n924), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n924), .B1(new_n941), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n934), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n910), .B1(new_n939), .B2(new_n940), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  INV_X1    g526(.A(new_n924), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n946), .A3(new_n933), .A4(new_n945), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n932), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n949), .C2(new_n954), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n947), .A2(new_n934), .A3(new_n948), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n957), .A2(new_n958), .B1(new_n959), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n510), .A2(new_n514), .B1(KEYINPUT4), .B2(new_n516), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n879), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT110), .B(G40), .Z(new_n969));
  NAND3_X1  g544(.A1(new_n473), .A2(new_n480), .A3(new_n969), .ZN(new_n970));
  OR3_X1    g545(.A1(new_n968), .A2(G1996), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n789), .B(G2067), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n803), .B2(G1996), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n968), .A2(new_n970), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n973), .A2(new_n803), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n733), .A2(new_n740), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G2067), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n875), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n976), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT127), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n973), .B(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n976), .B1(new_n974), .B2(new_n803), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n733), .A2(new_n740), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n976), .B1(new_n991), .B2(new_n980), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT48), .Z(new_n994));
  NAND3_X1  g569(.A1(new_n979), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n985), .A2(new_n986), .A3(new_n990), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n990), .A2(new_n995), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n977), .B1(new_n981), .B2(new_n983), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT127), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n979), .A2(new_n992), .ZN(new_n1001));
  XNOR2_X1  g576(.A(G290), .B(G1986), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n976), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n967), .A2(G1384), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n880), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT113), .B(new_n1005), .C1(new_n965), .C2(new_n879), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2078), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n468), .B1(new_n483), .B2(new_n484), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n469), .A2(new_n470), .ZN(new_n1012));
  OAI21_X1  g587(.A(G2105), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n472), .A2(G101), .ZN(new_n1014));
  AND4_X1   g589(.A1(new_n480), .A2(new_n1013), .A3(new_n1014), .A4(new_n969), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n967), .B1(G164), .B2(G1384), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(new_n1010), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n467), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n511), .B1(new_n478), .B2(new_n513), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n517), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n879), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n970), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n820), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1010), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1009), .A2(G160), .A3(new_n968), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1019), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1015), .B1(G164), .B2(new_n1006), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT53), .A3(new_n1010), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1019), .A2(new_n1037), .A3(new_n1029), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1033), .B(KEYINPUT54), .C1(G171), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1966), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT118), .B(G2084), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1026), .A2(new_n1027), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1043), .A3(G168), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  AOI21_X1  g620(.A(G168), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n506), .B1(new_n505), .B2(new_n493), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n505), .A2(new_n506), .A3(new_n493), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1022), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(new_n1025), .A3(new_n964), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT50), .B1(new_n880), .B2(G1384), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1015), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  AOI21_X1  g634(.A(G2090), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT117), .A4(new_n1015), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1060), .A2(new_n1061), .B1(new_n718), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1052), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1015), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1025), .B1(new_n1055), .B2(new_n964), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1062), .A2(new_n718), .B1(new_n1068), .B2(new_n761), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1069), .A2(new_n1064), .A3(new_n1052), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n704), .A2(G1976), .A3(new_n705), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1024), .A2(new_n1015), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(G8), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT114), .B(new_n1064), .C1(new_n1024), .C2(new_n1015), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1071), .B(new_n1073), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT115), .B(G86), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n601), .B(new_n603), .C1(new_n552), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G1981), .ZN(new_n1081));
  INV_X1    g656(.A(G1981), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n601), .A2(new_n1082), .A3(new_n602), .A4(new_n603), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1081), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT49), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n966), .A2(new_n970), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT114), .B1(new_n1088), .B2(new_n1064), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1075), .A2(new_n1074), .A3(G8), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1090), .B1(new_n707), .B2(G1976), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1078), .B(new_n1087), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1070), .A2(new_n1093), .ZN(new_n1094));
  AND4_X1   g669(.A1(new_n1039), .A2(new_n1050), .A3(new_n1065), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1038), .A2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT125), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1038), .A2(new_n1099), .A3(G171), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1032), .A2(G171), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .A4(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1015), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n815), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n577), .A2(new_n588), .A3(KEYINPUT57), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n525), .B1(new_n586), .B2(KEYINPUT78), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n583), .A2(new_n584), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1112), .A2(new_n1113), .B1(G91), .B2(new_n562), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n574), .A2(new_n576), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1106), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1109), .B2(new_n1106), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1117), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1106), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n970), .A2(G1996), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT113), .B1(new_n1131), .B2(new_n1005), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1008), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1016), .B(new_n1130), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1075), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1139), .A3(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1129), .B1(new_n1141), .B2(new_n565), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1134), .A2(new_n1139), .A3(new_n1136), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n565), .B(new_n1129), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1127), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1127), .B(new_n1149), .C1(new_n1142), .C2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n629), .A2(KEYINPUT123), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n623), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1088), .A2(new_n982), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1028), .A2(new_n810), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1155), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1152), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT123), .B(new_n629), .C1(new_n1158), .C2(new_n1152), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1148), .A2(new_n1150), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n623), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1118), .B1(new_n1163), .B2(new_n1123), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1104), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1078), .A2(new_n1087), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1092), .B1(new_n1168), .B2(new_n1071), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1052), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1062), .A2(new_n718), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1028), .A2(G2090), .ZN(new_n1173));
  OAI211_X1 g748(.A(G8), .B(new_n1171), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1064), .B(G286), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1065), .A2(new_n1170), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT119), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1052), .B1(new_n1069), .B2(new_n1064), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1094), .A2(new_n1182), .A3(KEYINPUT63), .A4(new_n1175), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n596), .A2(new_n1072), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT116), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1083), .B1(new_n1186), .B2(new_n1086), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1168), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1174), .B2(new_n1093), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1065), .A2(new_n1174), .A3(new_n1170), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n1100), .B2(new_n1098), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1047), .A2(new_n1192), .A3(new_n1049), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1189), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1184), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT126), .B(new_n1003), .C1(new_n1166), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1161), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1147), .B2(KEYINPUT122), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1164), .B1(new_n1201), .B2(new_n1150), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1184), .B(new_n1196), .C1(new_n1202), .C2(new_n1104), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT126), .B1(new_n1203), .B2(new_n1003), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1000), .B1(new_n1199), .B2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g780(.A1(G229), .A2(G227), .A3(new_n463), .A4(G401), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n896), .A2(new_n955), .A3(new_n1207), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


