

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n902), .Z(n513) );
  XOR2_X1 U551 ( .A(n648), .B(KEYINPUT15), .Z(n984) );
  NOR2_X1 U552 ( .A1(n549), .A2(n548), .ZN(G164) );
  NOR2_X4 U553 ( .A1(n618), .A2(n617), .ZN(G160) );
  XNOR2_X1 U554 ( .A(n541), .B(n540), .ZN(n902) );
  NOR2_X1 U555 ( .A1(n690), .A2(n689), .ZN(n692) );
  AND2_X1 U556 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U557 ( .A(n697), .B(KEYINPUT30), .ZN(n698) );
  OR2_X1 U558 ( .A1(n717), .A2(n696), .ZN(n697) );
  OR2_X1 U559 ( .A1(n719), .A2(n695), .ZN(n696) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n625) );
  BUF_X2 U561 ( .A(n794), .Z(n514) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n519), .Z(n794) );
  XNOR2_X1 U563 ( .A(n638), .B(KEYINPUT28), .ZN(n676) );
  XNOR2_X1 U564 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n701) );
  AND2_X1 U565 ( .A1(n518), .A2(n973), .ZN(n736) );
  NOR2_X1 U566 ( .A1(G543), .A2(n525), .ZN(n519) );
  XNOR2_X2 U567 ( .A(n543), .B(KEYINPUT65), .ZN(n579) );
  AND2_X1 U568 ( .A1(n546), .A2(n545), .ZN(n515) );
  OR2_X1 U569 ( .A1(n745), .A2(n744), .ZN(n516) );
  AND2_X1 U570 ( .A1(n746), .A2(n516), .ZN(n517) );
  OR2_X1 U571 ( .A1(n735), .A2(n745), .ZN(n518) );
  BUF_X1 U572 ( .A(n694), .Z(n703) );
  INV_X1 U573 ( .A(KEYINPUT100), .ZN(n691) );
  XNOR2_X1 U574 ( .A(n702), .B(n701), .ZN(n716) );
  INV_X1 U575 ( .A(KEYINPUT103), .ZN(n729) );
  INV_X1 U576 ( .A(n686), .ZN(n694) );
  INV_X1 U577 ( .A(KEYINPUT17), .ZN(n540) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n541) );
  NOR2_X2 U579 ( .A1(G2105), .A2(n544), .ZN(n901) );
  NOR2_X1 U580 ( .A1(G651), .A2(n565), .ZN(n793) );
  XNOR2_X1 U581 ( .A(n758), .B(KEYINPUT40), .ZN(n759) );
  XOR2_X1 U582 ( .A(G651), .B(KEYINPUT66), .Z(n525) );
  NAND2_X1 U583 ( .A1(G63), .A2(n514), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT74), .ZN(n522) );
  XOR2_X1 U585 ( .A(G543), .B(KEYINPUT0), .Z(n565) );
  NAND2_X1 U586 ( .A1(G51), .A2(n793), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n523), .ZN(n530) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n799) );
  NAND2_X1 U590 ( .A1(n799), .A2(G89), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n565), .A2(n525), .ZN(n797) );
  NAND2_X1 U593 ( .A1(G76), .A2(n797), .ZN(n526) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U595 ( .A(n528), .B(KEYINPUT5), .Z(n529) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT7), .B(n531), .Z(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT75), .B(n532), .Z(G168) );
  NAND2_X1 U599 ( .A1(n799), .A2(G85), .ZN(n534) );
  NAND2_X1 U600 ( .A1(G72), .A2(n797), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U602 ( .A1(G47), .A2(n793), .ZN(n535) );
  XNOR2_X1 U603 ( .A(KEYINPUT67), .B(n535), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U605 ( .A1(G60), .A2(n514), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(G290) );
  NAND2_X1 U607 ( .A1(n902), .A2(G138), .ZN(n542) );
  XOR2_X1 U608 ( .A(n542), .B(KEYINPUT90), .Z(n549) );
  INV_X1 U609 ( .A(G2104), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n544), .A2(G2105), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n579), .A2(G126), .ZN(n547) );
  AND2_X1 U612 ( .A1(G2105), .A2(G2104), .ZN(n905) );
  NAND2_X1 U613 ( .A1(G114), .A2(n905), .ZN(n546) );
  NAND2_X1 U614 ( .A1(G102), .A2(n901), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n547), .A2(n515), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n799), .A2(G90), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G77), .A2(n797), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT69), .B(KEYINPUT9), .Z(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n514), .A2(G64), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n793), .A2(G52), .ZN(n555) );
  AND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(G301) );
  NAND2_X1 U626 ( .A1(n799), .A2(G88), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G75), .A2(n797), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n793), .A2(G50), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G62), .A2(n514), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U632 ( .A1(n564), .A2(n563), .ZN(G166) );
  INV_X1 U633 ( .A(G166), .ZN(G303) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G87), .A2(n565), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U638 ( .A1(n514), .A2(n568), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n793), .A2(G49), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U641 ( .A1(n799), .A2(G86), .ZN(n572) );
  NAND2_X1 U642 ( .A1(G61), .A2(n514), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U644 ( .A(KEYINPUT84), .B(n573), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G73), .A2(n797), .ZN(n574) );
  XOR2_X1 U646 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n793), .A2(G48), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U650 ( .A1(G117), .A2(n905), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G129), .A2(n579), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n901), .A2(G105), .ZN(n582) );
  XOR2_X1 U654 ( .A(KEYINPUT38), .B(n582), .Z(n583) );
  NOR2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n513), .A2(G141), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n883) );
  NOR2_X1 U658 ( .A1(G1996), .A2(n883), .ZN(n935) );
  NAND2_X1 U659 ( .A1(G107), .A2(n905), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G119), .A2(n579), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n901), .A2(G95), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT92), .B(n589), .Z(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n513), .A2(G131), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n897) );
  NAND2_X1 U667 ( .A1(G1991), .A2(n897), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT93), .B(n594), .Z(n596) );
  NAND2_X1 U669 ( .A1(G1996), .A2(n883), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n925) );
  NOR2_X1 U671 ( .A1(G1986), .A2(G290), .ZN(n597) );
  NOR2_X1 U672 ( .A1(G1991), .A2(n897), .ZN(n926) );
  NOR2_X1 U673 ( .A1(n597), .A2(n926), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT105), .B(n598), .Z(n599) );
  NOR2_X1 U675 ( .A1(n925), .A2(n599), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n935), .A2(n600), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT39), .ZN(n619) );
  NAND2_X1 U678 ( .A1(G104), .A2(n901), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G140), .A2(n513), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT91), .B(KEYINPUT34), .Z(n604) );
  XNOR2_X1 U682 ( .A(n605), .B(n604), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G116), .A2(n905), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G128), .A2(n579), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT35), .B(n608), .Z(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U688 ( .A(KEYINPUT36), .B(n611), .ZN(n887) );
  INV_X1 U689 ( .A(G2067), .ZN(n855) );
  XOR2_X1 U690 ( .A(KEYINPUT37), .B(n855), .Z(n620) );
  NOR2_X1 U691 ( .A1(n887), .A2(n620), .ZN(n943) );
  NAND2_X1 U692 ( .A1(n905), .A2(G113), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G101), .A2(n901), .ZN(n612) );
  XOR2_X1 U694 ( .A(KEYINPUT23), .B(n612), .Z(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G125), .A2(n579), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G137), .A2(n513), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U699 ( .A1(G160), .A2(G40), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n625), .A2(n626), .ZN(n749) );
  NAND2_X1 U701 ( .A1(n943), .A2(n749), .ZN(n753) );
  NAND2_X1 U702 ( .A1(n619), .A2(n753), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n887), .A2(n620), .ZN(n941) );
  NAND2_X1 U704 ( .A1(n621), .A2(n941), .ZN(n622) );
  XNOR2_X1 U705 ( .A(KEYINPUT106), .B(n622), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n623), .A2(n749), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n624), .B(KEYINPUT107), .ZN(n757) );
  INV_X1 U708 ( .A(n625), .ZN(n627) );
  NOR2_X2 U709 ( .A1(n627), .A2(n626), .ZN(n686) );
  NAND2_X1 U710 ( .A1(n686), .A2(G2072), .ZN(n628) );
  XNOR2_X1 U711 ( .A(n628), .B(KEYINPUT27), .ZN(n630) );
  INV_X1 U712 ( .A(G1956), .ZN(n866) );
  NOR2_X1 U713 ( .A1(n866), .A2(n686), .ZN(n629) );
  NOR2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n799), .A2(G91), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G78), .A2(n797), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n793), .A2(G53), .ZN(n634) );
  NAND2_X1 U719 ( .A1(G65), .A2(n514), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U722 ( .A(KEYINPUT70), .B(n637), .ZN(n989) );
  NOR2_X1 U723 ( .A1(n639), .A2(n989), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n639), .A2(n989), .ZN(n640) );
  OR2_X1 U725 ( .A1(n676), .A2(n640), .ZN(n683) );
  NAND2_X1 U726 ( .A1(G54), .A2(n793), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n799), .A2(G92), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G66), .A2(n514), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U730 ( .A1(G79), .A2(n797), .ZN(n643) );
  XNOR2_X1 U731 ( .A(KEYINPUT73), .B(n643), .ZN(n644) );
  NOR2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n648) );
  INV_X1 U734 ( .A(n984), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G1348), .A2(n694), .ZN(n649) );
  XNOR2_X1 U736 ( .A(KEYINPUT98), .B(n649), .ZN(n651) );
  NOR2_X1 U737 ( .A1(n855), .A2(n694), .ZN(n650) );
  NAND2_X1 U738 ( .A1(KEYINPUT98), .A2(n650), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n651), .A2(n654), .ZN(n653) );
  INV_X1 U740 ( .A(KEYINPUT99), .ZN(n652) );
  NAND2_X1 U741 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U742 ( .A1(n654), .A2(KEYINPUT99), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n656), .A2(n655), .ZN(n677) );
  INV_X1 U744 ( .A(n677), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n658), .A2(n657), .ZN(n675) );
  INV_X1 U746 ( .A(G1996), .ZN(n867) );
  NOR2_X1 U747 ( .A1(n694), .A2(n867), .ZN(n660) );
  XOR2_X1 U748 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n659) );
  XNOR2_X1 U749 ( .A(n660), .B(n659), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n703), .A2(G1341), .ZN(n661) );
  NAND2_X1 U751 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U752 ( .A(KEYINPUT97), .B(n663), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n799), .A2(G81), .ZN(n664) );
  XNOR2_X1 U754 ( .A(n664), .B(KEYINPUT12), .ZN(n666) );
  NAND2_X1 U755 ( .A1(G68), .A2(n797), .ZN(n665) );
  NAND2_X1 U756 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U757 ( .A(n667), .B(KEYINPUT13), .ZN(n669) );
  NAND2_X1 U758 ( .A1(G43), .A2(n793), .ZN(n668) );
  NAND2_X1 U759 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n514), .A2(G56), .ZN(n670) );
  XOR2_X1 U761 ( .A(KEYINPUT14), .B(n670), .Z(n671) );
  NOR2_X1 U762 ( .A1(n672), .A2(n671), .ZN(n988) );
  NAND2_X1 U763 ( .A1(n673), .A2(n988), .ZN(n674) );
  NAND2_X1 U764 ( .A1(n675), .A2(n674), .ZN(n681) );
  INV_X1 U765 ( .A(n676), .ZN(n679) );
  NAND2_X1 U766 ( .A1(n984), .A2(n677), .ZN(n678) );
  AND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n684), .B(KEYINPUT29), .ZN(n690) );
  NAND2_X1 U770 ( .A1(G1961), .A2(n703), .ZN(n688) );
  XOR2_X1 U771 ( .A(G2078), .B(KEYINPUT96), .Z(n685) );
  XNOR2_X1 U772 ( .A(KEYINPUT25), .B(n685), .ZN(n951) );
  NAND2_X1 U773 ( .A1(n686), .A2(n951), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n693) );
  NOR2_X1 U775 ( .A1(G301), .A2(n693), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n692), .B(n691), .ZN(n715) );
  AND2_X1 U777 ( .A1(G301), .A2(n693), .ZN(n700) );
  NAND2_X1 U778 ( .A1(G8), .A2(n694), .ZN(n745) );
  NOR2_X1 U779 ( .A1(G1966), .A2(n745), .ZN(n717) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n703), .ZN(n719) );
  INV_X1 U781 ( .A(G8), .ZN(n695) );
  NOR2_X1 U782 ( .A1(n698), .A2(G168), .ZN(n699) );
  NOR2_X1 U783 ( .A1(n700), .A2(n699), .ZN(n702) );
  NOR2_X1 U784 ( .A1(G1971), .A2(n745), .ZN(n705) );
  NOR2_X1 U785 ( .A1(G2090), .A2(n703), .ZN(n704) );
  NOR2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U787 ( .A1(n706), .A2(G303), .ZN(n707) );
  OR2_X1 U788 ( .A1(n695), .A2(n707), .ZN(n709) );
  AND2_X1 U789 ( .A1(n716), .A2(n709), .ZN(n708) );
  NAND2_X1 U790 ( .A1(n715), .A2(n708), .ZN(n713) );
  INV_X1 U791 ( .A(n709), .ZN(n711) );
  AND2_X1 U792 ( .A1(G286), .A2(G8), .ZN(n710) );
  OR2_X1 U793 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U795 ( .A(n714), .B(KEYINPUT32), .ZN(n724) );
  AND2_X1 U796 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U797 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U798 ( .A1(G8), .A2(n719), .ZN(n720) );
  XOR2_X1 U799 ( .A(KEYINPUT95), .B(n720), .Z(n721) );
  NAND2_X1 U800 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U801 ( .A1(n724), .A2(n723), .ZN(n739) );
  NOR2_X1 U802 ( .A1(G1971), .A2(G303), .ZN(n725) );
  XOR2_X1 U803 ( .A(n725), .B(KEYINPUT102), .Z(n726) );
  NOR2_X1 U804 ( .A1(G1976), .A2(G288), .ZN(n734) );
  INV_X1 U805 ( .A(n734), .ZN(n977) );
  AND2_X1 U806 ( .A1(n726), .A2(n977), .ZN(n727) );
  NAND2_X1 U807 ( .A1(n739), .A2(n727), .ZN(n728) );
  NAND2_X1 U808 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NAND2_X1 U809 ( .A1(n728), .A2(n976), .ZN(n730) );
  XNOR2_X1 U810 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U811 ( .A1(n731), .A2(n745), .ZN(n732) );
  NOR2_X1 U812 ( .A1(KEYINPUT33), .A2(n732), .ZN(n733) );
  INV_X1 U813 ( .A(n733), .ZN(n737) );
  NAND2_X1 U814 ( .A1(n734), .A2(KEYINPUT33), .ZN(n735) );
  XOR2_X1 U815 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U816 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U817 ( .A(n738), .B(KEYINPUT104), .ZN(n747) );
  NOR2_X1 U818 ( .A1(G2090), .A2(G303), .ZN(n740) );
  NAND2_X1 U819 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U820 ( .A1(n739), .A2(n741), .ZN(n742) );
  NAND2_X1 U821 ( .A1(n742), .A2(n745), .ZN(n746) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n743) );
  XOR2_X1 U823 ( .A(n743), .B(KEYINPUT24), .Z(n744) );
  AND2_X1 U824 ( .A1(n747), .A2(n517), .ZN(n755) );
  NAND2_X1 U825 ( .A1(n925), .A2(n749), .ZN(n748) );
  XNOR2_X1 U826 ( .A(n748), .B(KEYINPUT94), .ZN(n751) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U828 ( .A1(n980), .A2(n749), .ZN(n750) );
  AND2_X1 U829 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n760) );
  INV_X1 U833 ( .A(KEYINPUT108), .ZN(n758) );
  XNOR2_X1 U834 ( .A(n760), .B(n759), .ZN(G329) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n764) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n762) );
  XOR2_X1 U840 ( .A(n762), .B(KEYINPUT10), .Z(n922) );
  NAND2_X1 U841 ( .A1(G567), .A2(n922), .ZN(n763) );
  XNOR2_X1 U842 ( .A(n764), .B(n763), .ZN(G234) );
  NAND2_X1 U843 ( .A1(n988), .A2(G860), .ZN(G153) );
  NAND2_X1 U844 ( .A1(G868), .A2(G301), .ZN(n766) );
  INV_X1 U845 ( .A(G868), .ZN(n810) );
  NAND2_X1 U846 ( .A1(n984), .A2(n810), .ZN(n765) );
  NAND2_X1 U847 ( .A1(n766), .A2(n765), .ZN(G284) );
  INV_X1 U848 ( .A(n989), .ZN(G299) );
  NOR2_X1 U849 ( .A1(G286), .A2(n810), .ZN(n768) );
  NOR2_X1 U850 ( .A1(G299), .A2(G868), .ZN(n767) );
  NOR2_X1 U851 ( .A1(n768), .A2(n767), .ZN(G297) );
  INV_X1 U852 ( .A(G860), .ZN(n843) );
  NAND2_X1 U853 ( .A1(G559), .A2(n843), .ZN(n769) );
  XOR2_X1 U854 ( .A(KEYINPUT76), .B(n769), .Z(n770) );
  NOR2_X1 U855 ( .A1(n984), .A2(n770), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT77), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U858 ( .A1(n988), .A2(n810), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT78), .B(n773), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n984), .A2(G559), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G868), .A2(n774), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U863 ( .A(KEYINPUT79), .B(n777), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G111), .A2(n905), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G99), .A2(n901), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT80), .B(n780), .ZN(n785) );
  NAND2_X1 U868 ( .A1(n579), .A2(G123), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G135), .A2(n513), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n924) );
  XNOR2_X1 U873 ( .A(n924), .B(G2096), .ZN(n786) );
  INV_X1 U874 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U875 ( .A1(n786), .A2(n852), .ZN(G156) );
  XNOR2_X1 U876 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n788) );
  XNOR2_X1 U877 ( .A(G288), .B(KEYINPUT19), .ZN(n787) );
  XNOR2_X1 U878 ( .A(n788), .B(n787), .ZN(n789) );
  XNOR2_X1 U879 ( .A(G290), .B(n789), .ZN(n791) );
  XOR2_X1 U880 ( .A(n989), .B(G166), .Z(n790) );
  XNOR2_X1 U881 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(G305), .ZN(n806) );
  NAND2_X1 U883 ( .A1(n793), .A2(G55), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G67), .A2(n514), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n798) );
  XOR2_X1 U887 ( .A(KEYINPUT81), .B(n798), .Z(n801) );
  NAND2_X1 U888 ( .A1(n799), .A2(G93), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(KEYINPUT82), .B(n802), .ZN(n803) );
  NOR2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n805), .B(KEYINPUT83), .ZN(n844) );
  XNOR2_X1 U893 ( .A(n806), .B(n844), .ZN(n846) );
  NAND2_X1 U894 ( .A1(G559), .A2(n658), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(n988), .ZN(n842) );
  XNOR2_X1 U896 ( .A(n846), .B(n842), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n808), .A2(G868), .ZN(n809) );
  XOR2_X1 U898 ( .A(KEYINPUT87), .B(n809), .Z(n812) );
  NAND2_X1 U899 ( .A1(n844), .A2(n810), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U907 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n817) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n817), .Z(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT88), .ZN(n819) );
  NOR2_X1 U911 ( .A1(G218), .A2(n819), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G96), .A2(n820), .ZN(n840) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n840), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G120), .A2(G69), .ZN(n821) );
  NOR2_X1 U915 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G108), .A2(n822), .ZN(n841) );
  NAND2_X1 U917 ( .A1(G567), .A2(n841), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U919 ( .A(KEYINPUT89), .B(n825), .Z(n851) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n851), .A2(n826), .ZN(n839) );
  NAND2_X1 U922 ( .A1(n839), .A2(G36), .ZN(G176) );
  XOR2_X1 U923 ( .A(G2430), .B(G2451), .Z(n828) );
  XNOR2_X1 U924 ( .A(G2446), .B(G2427), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(n835) );
  XOR2_X1 U926 ( .A(G2438), .B(G2435), .Z(n830) );
  XNOR2_X1 U927 ( .A(G2443), .B(KEYINPUT109), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U929 ( .A(n831), .B(G2454), .Z(n833) );
  XNOR2_X1 U930 ( .A(G1348), .B(G1341), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n836), .A2(G14), .ZN(n915) );
  XOR2_X1 U934 ( .A(KEYINPUT110), .B(n915), .Z(G401) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n922), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U937 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U939 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U940 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n841), .A2(n840), .ZN(G325) );
  XOR2_X1 U942 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  NAND2_X1 U945 ( .A1(n843), .A2(n842), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(G145) );
  XOR2_X1 U947 ( .A(n846), .B(G286), .Z(n848) );
  XOR2_X1 U948 ( .A(G301), .B(n988), .Z(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n849), .B(n984), .Z(n850) );
  NOR2_X1 U951 ( .A1(G37), .A2(n850), .ZN(G397) );
  INV_X1 U952 ( .A(n851), .ZN(G319) );
  XNOR2_X1 U953 ( .A(n852), .B(G2096), .ZN(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n859) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XOR2_X1 U957 ( .A(n855), .B(G2072), .Z(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1976), .B(G1981), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1971), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n875) );
  XOR2_X1 U965 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n865) );
  XNOR2_X1 U966 ( .A(G1991), .B(KEYINPUT41), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n871) );
  XNOR2_X1 U968 ( .A(G1986), .B(n866), .ZN(n869) );
  XOR2_X1 U969 ( .A(G1961), .B(n867), .Z(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT113), .B(G2474), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(n875), .B(n874), .Z(G229) );
  NAND2_X1 U975 ( .A1(G112), .A2(n905), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G100), .A2(n901), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U978 ( .A1(n579), .A2(G124), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G136), .A2(n513), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(G162) );
  XNOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n883), .B(n924), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(G162), .B(n886), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n887), .B(G164), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n900) );
  NAND2_X1 U989 ( .A1(G118), .A2(n905), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G130), .A2(n579), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G106), .A2(n901), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G142), .A2(n513), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(n894), .B(KEYINPUT45), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n913) );
  NAND2_X1 U999 ( .A1(G103), .A2(n901), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G139), .A2(n513), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n905), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n579), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT116), .B(n911), .Z(n929) );
  XNOR2_X1 U1008 ( .A(G160), .B(n929), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G397), .A2(n916), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n920), .A2(G395), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n921), .B(KEYINPUT117), .Z(G308) );
  INV_X1 U1018 ( .A(G308), .ZN(G225) );
  INV_X1 U1019 ( .A(G96), .ZN(G221) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  INV_X1 U1021 ( .A(n922), .ZN(G223) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n940) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n931) );
  XNOR2_X1 U1027 ( .A(G2072), .B(n929), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n932), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT50), .ZN(n938) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n945) );
  INV_X1 U1036 ( .A(n941), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(n947), .ZN(n948) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n968) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n968), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n949), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1044 ( .A(G29), .B(KEYINPUT122), .Z(n971) );
  XOR2_X1 U1045 ( .A(G2090), .B(G35), .Z(n964) );
  XOR2_X1 U1046 ( .A(G2072), .B(G33), .Z(n950) );
  NAND2_X1 U1047 ( .A1(n950), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G27), .B(n951), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(KEYINPUT120), .B(n952), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1051 ( .A(G1996), .B(G32), .Z(n956) );
  XOR2_X1 U1052 ( .A(G2067), .B(G26), .Z(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT121), .B(n961), .Z(n962) );
  XNOR2_X1 U1058 ( .A(n962), .B(KEYINPUT53), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G34), .B(G2084), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n969), .B(n968), .Z(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n972), .ZN(n1027) );
  INV_X1 U1066 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1067 ( .A(n1023), .B(KEYINPUT56), .Z(n999) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(KEYINPUT57), .ZN(n997) );
  XOR2_X1 U1071 ( .A(G303), .B(G1971), .Z(n982) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT125), .B(n978), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n995) );
  XOR2_X1 U1076 ( .A(G301), .B(G1961), .Z(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G1348), .B(n984), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n987), .ZN(n993) );
  XOR2_X1 U1081 ( .A(n988), .B(G1341), .Z(n991) );
  XOR2_X1 U1082 ( .A(n989), .B(G1956), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1025) );
  XOR2_X1 U1088 ( .A(G20), .B(G1956), .Z(n1003) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G6), .B(G1981), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1007), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1008), .B(KEYINPUT126), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G5), .B(G1961), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT61), .Z(n1021) );
  XNOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
  INV_X1 U1117 ( .A(G301), .ZN(G171) );
endmodule

