

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601;

  NOR2_X1 U325 ( .A1(n553), .A2(n468), .ZN(n573) );
  XNOR2_X1 U326 ( .A(n332), .B(n331), .ZN(n335) );
  XNOR2_X1 U327 ( .A(n398), .B(n397), .ZN(n523) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n422) );
  XNOR2_X1 U329 ( .A(n467), .B(n466), .ZN(n577) );
  NOR2_X1 U330 ( .A1(n553), .A2(n499), .ZN(n589) );
  XOR2_X1 U331 ( .A(n372), .B(n371), .Z(n293) );
  XOR2_X1 U332 ( .A(n418), .B(KEYINPUT114), .Z(n294) );
  NOR2_X1 U333 ( .A1(n578), .A2(n530), .ZN(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT106), .B(n487), .Z(n296) );
  XOR2_X1 U335 ( .A(n409), .B(n408), .Z(n297) );
  XOR2_X1 U336 ( .A(G99GAT), .B(G85GAT), .Z(n376) );
  XNOR2_X1 U337 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U338 ( .A(n384), .B(n383), .ZN(n385) );
  INV_X1 U339 ( .A(KEYINPUT92), .ZN(n329) );
  XNOR2_X1 U340 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U341 ( .A(n386), .B(n385), .ZN(n389) );
  XNOR2_X1 U342 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U343 ( .A(KEYINPUT37), .B(KEYINPUT107), .ZN(n488) );
  XNOR2_X1 U344 ( .A(n373), .B(n293), .ZN(n374) );
  INV_X1 U345 ( .A(KEYINPUT116), .ZN(n466) );
  XNOR2_X1 U346 ( .A(n489), .B(n488), .ZN(n510) );
  XNOR2_X1 U347 ( .A(n375), .B(n374), .ZN(n508) );
  XNOR2_X1 U348 ( .A(n591), .B(n422), .ZN(n500) );
  XNOR2_X1 U349 ( .A(n518), .B(KEYINPUT125), .ZN(n519) );
  XOR2_X1 U350 ( .A(n415), .B(n414), .Z(n595) );
  XNOR2_X1 U351 ( .A(n490), .B(KEYINPUT111), .ZN(n565) );
  XNOR2_X1 U352 ( .A(n520), .B(n519), .ZN(n522) );
  XNOR2_X1 U353 ( .A(n469), .B(G127GAT), .ZN(n470) );
  XNOR2_X1 U354 ( .A(KEYINPUT112), .B(G85GAT), .ZN(n491) );
  XNOR2_X1 U355 ( .A(n507), .B(n506), .ZN(G1351GAT) );
  XNOR2_X1 U356 ( .A(n492), .B(n491), .ZN(G1336GAT) );
  XNOR2_X1 U357 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n298), .B(KEYINPUT17), .ZN(n299) );
  XOR2_X1 U359 ( .A(n299), .B(KEYINPUT18), .Z(n301) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(G176GAT), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n433) );
  XOR2_X1 U362 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT84), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n460) );
  XNOR2_X1 U365 ( .A(n460), .B(KEYINPUT20), .ZN(n304) );
  AND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  NAND2_X1 U367 ( .A1(n304), .A2(n305), .ZN(n309) );
  INV_X1 U368 ( .A(n304), .ZN(n307) );
  INV_X1 U369 ( .A(n305), .ZN(n306) );
  NAND2_X1 U370 ( .A1(n307), .A2(n306), .ZN(n308) );
  NAND2_X1 U371 ( .A1(n309), .A2(n308), .ZN(n310) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G71GAT), .Z(n357) );
  XNOR2_X1 U373 ( .A(n310), .B(n357), .ZN(n312) );
  XOR2_X1 U374 ( .A(G99GAT), .B(G190GAT), .Z(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n314) );
  XOR2_X1 U376 ( .A(G43GAT), .B(G134GAT), .Z(n382) );
  XOR2_X1 U377 ( .A(G15GAT), .B(G127GAT), .Z(n402) );
  XNOR2_X1 U378 ( .A(n382), .B(n402), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U380 ( .A(n433), .B(n315), .Z(n472) );
  INV_X1 U381 ( .A(n472), .ZN(n553) );
  XOR2_X1 U382 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n317) );
  XNOR2_X1 U383 ( .A(KEYINPUT90), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U384 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U385 ( .A(KEYINPUT3), .B(n318), .ZN(n455) );
  XOR2_X1 U386 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n320) );
  XNOR2_X1 U387 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n319) );
  XNOR2_X1 U388 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U389 ( .A(n455), .B(n321), .Z(n337) );
  INV_X1 U390 ( .A(G197GAT), .ZN(n325) );
  XOR2_X1 U391 ( .A(KEYINPUT89), .B(G218GAT), .Z(n323) );
  XNOR2_X1 U392 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U393 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n325), .B(n324), .ZN(n432) );
  XOR2_X1 U395 ( .A(KEYINPUT22), .B(G204GAT), .Z(n327) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n344) );
  XOR2_X1 U397 ( .A(G50GAT), .B(G162GAT), .Z(n377) );
  XNOR2_X1 U398 ( .A(n344), .B(n377), .ZN(n326) );
  XNOR2_X1 U399 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U400 ( .A(n432), .B(n328), .Z(n332) );
  NAND2_X1 U401 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U403 ( .A(n333), .B(G148GAT), .ZN(n364) );
  XNOR2_X1 U404 ( .A(n364), .B(KEYINPUT87), .ZN(n334) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n497) );
  XNOR2_X1 U407 ( .A(n497), .B(KEYINPUT28), .ZN(n564) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G113GAT), .Z(n339) );
  XNOR2_X1 U409 ( .A(G43GAT), .B(G50GAT), .ZN(n338) );
  XNOR2_X1 U410 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U411 ( .A(n340), .B(G36GAT), .Z(n342) );
  XOR2_X1 U412 ( .A(G1GAT), .B(G8GAT), .Z(n403) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(n403), .ZN(n341) );
  XNOR2_X1 U414 ( .A(n342), .B(n341), .ZN(n348) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n343) );
  XNOR2_X1 U416 ( .A(n343), .B(KEYINPUT8), .ZN(n396) );
  XOR2_X1 U417 ( .A(n396), .B(n344), .Z(n346) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U420 ( .A(n348), .B(n347), .Z(n356) );
  XOR2_X1 U421 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n350) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(KEYINPUT69), .ZN(n349) );
  XNOR2_X1 U423 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U424 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n352) );
  XNOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n351) );
  XNOR2_X1 U426 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n356), .B(n355), .ZN(n587) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n359) );
  XNOR2_X1 U430 ( .A(n357), .B(n376), .ZN(n358) );
  XNOR2_X1 U431 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U432 ( .A(n360), .B(KEYINPUT32), .Z(n367) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  INV_X1 U434 ( .A(KEYINPUT72), .ZN(n361) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n375) );
  XNOR2_X1 U437 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n368), .B(KEYINPUT13), .ZN(n404) );
  XOR2_X1 U439 ( .A(G64GAT), .B(KEYINPUT74), .Z(n370) );
  XNOR2_X1 U440 ( .A(G204GAT), .B(G92GAT), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n436) );
  XNOR2_X1 U442 ( .A(n404), .B(n436), .ZN(n373) );
  XOR2_X1 U443 ( .A(KEYINPUT76), .B(KEYINPUT73), .Z(n372) );
  XNOR2_X1 U444 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n371) );
  INV_X1 U445 ( .A(n508), .ZN(n591) );
  XOR2_X1 U446 ( .A(KEYINPUT9), .B(n376), .Z(n379) );
  XNOR2_X1 U447 ( .A(G218GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n386) );
  XOR2_X1 U449 ( .A(G92GAT), .B(KEYINPUT81), .Z(n381) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n380) );
  XOR2_X1 U451 ( .A(n381), .B(n380), .Z(n384) );
  XNOR2_X1 U452 ( .A(n382), .B(KEYINPUT10), .ZN(n383) );
  XOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n388) );
  XNOR2_X1 U454 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n387) );
  XOR2_X1 U455 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U456 ( .A1(n389), .A2(n390), .ZN(n394) );
  INV_X1 U457 ( .A(n389), .ZN(n392) );
  INV_X1 U458 ( .A(n390), .ZN(n391) );
  NAND2_X1 U459 ( .A1(n392), .A2(n391), .ZN(n393) );
  NAND2_X1 U460 ( .A1(n394), .A2(n393), .ZN(n398) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(G190GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n395), .B(KEYINPUT80), .ZN(n438) );
  XOR2_X1 U463 ( .A(n396), .B(n438), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n399) );
  XOR2_X1 U465 ( .A(n523), .B(n399), .Z(n599) );
  XOR2_X1 U466 ( .A(G155GAT), .B(G78GAT), .Z(n401) );
  XNOR2_X1 U467 ( .A(G183GAT), .B(G71GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U471 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n407) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U474 ( .A(KEYINPUT82), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U475 ( .A(G22GAT), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n412), .B(KEYINPUT15), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n297), .B(n413), .ZN(n414) );
  INV_X1 U479 ( .A(n595), .ZN(n421) );
  NOR2_X1 U480 ( .A1(n599), .A2(n421), .ZN(n416) );
  XOR2_X1 U481 ( .A(n416), .B(KEYINPUT45), .Z(n417) );
  NOR2_X1 U482 ( .A1(n591), .A2(n417), .ZN(n418) );
  OR2_X1 U483 ( .A1(n587), .A2(n294), .ZN(n420) );
  INV_X1 U484 ( .A(KEYINPUT115), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n430) );
  NAND2_X1 U486 ( .A1(n523), .A2(n421), .ZN(n427) );
  XNOR2_X1 U487 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n425) );
  INV_X1 U488 ( .A(n500), .ZN(n423) );
  NAND2_X1 U489 ( .A1(n587), .A2(n423), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U491 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(KEYINPUT47), .B(n428), .ZN(n429) );
  AND2_X1 U493 ( .A1(n430), .A2(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n431), .B(KEYINPUT48), .ZN(n494) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n442) );
  XOR2_X1 U496 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n435) );
  NAND2_X1 U497 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U499 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U500 ( .A(G8GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(n441), .Z(n551) );
  XNOR2_X1 U503 ( .A(n551), .B(KEYINPUT27), .ZN(n477) );
  XOR2_X1 U504 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n444) );
  XNOR2_X1 U505 ( .A(G141GAT), .B(G148GAT), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U507 ( .A(G85GAT), .B(G120GAT), .Z(n446) );
  XNOR2_X1 U508 ( .A(G29GAT), .B(G127GAT), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n450) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n452) );
  XNOR2_X1 U515 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U520 ( .A(G134GAT), .B(n459), .ZN(n464) );
  XOR2_X1 U521 ( .A(G162GAT), .B(n460), .Z(n462) );
  NAND2_X1 U522 ( .A1(G225GAT), .A2(G233GAT), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U524 ( .A(n464), .B(n463), .Z(n530) );
  INV_X1 U525 ( .A(n530), .ZN(n548) );
  NOR2_X1 U526 ( .A1(n477), .A2(n548), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT100), .B(n465), .Z(n483) );
  NOR2_X1 U528 ( .A1(n494), .A2(n483), .ZN(n467) );
  OR2_X1 U529 ( .A1(n564), .A2(n577), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n573), .A2(n595), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n469) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(G1342GAT) );
  NOR2_X1 U533 ( .A1(n587), .A2(n500), .ZN(n547) );
  INV_X1 U534 ( .A(n551), .ZN(n560) );
  NAND2_X1 U535 ( .A1(n472), .A2(n560), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n473), .B(KEYINPUT101), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n474), .A2(n497), .ZN(n475) );
  XOR2_X1 U538 ( .A(KEYINPUT25), .B(n475), .Z(n479) );
  NAND2_X1 U539 ( .A1(n553), .A2(n497), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n476), .B(KEYINPUT26), .ZN(n578) );
  NOR2_X1 U541 ( .A1(n578), .A2(n477), .ZN(n478) );
  NOR2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U543 ( .A1(n480), .A2(n530), .ZN(n485) );
  INV_X1 U544 ( .A(n553), .ZN(n562) );
  XOR2_X1 U545 ( .A(KEYINPUT86), .B(n562), .Z(n481) );
  INV_X1 U546 ( .A(n564), .ZN(n556) );
  NAND2_X1 U547 ( .A1(n481), .A2(n556), .ZN(n482) );
  NOR2_X1 U548 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U549 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n486), .B(KEYINPUT102), .ZN(n526) );
  NOR2_X1 U551 ( .A1(n595), .A2(n526), .ZN(n487) );
  NOR2_X1 U552 ( .A1(n599), .A2(n296), .ZN(n489) );
  NAND2_X1 U553 ( .A1(n547), .A2(n510), .ZN(n490) );
  NAND2_X1 U554 ( .A1(n530), .A2(n565), .ZN(n492) );
  XOR2_X1 U555 ( .A(n551), .B(KEYINPUT121), .Z(n493) );
  NOR2_X1 U556 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT54), .ZN(n516) );
  NAND2_X1 U558 ( .A1(n516), .A2(n548), .ZN(n496) );
  NOR2_X1 U559 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT55), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n589), .A2(n423), .ZN(n503) );
  XOR2_X1 U562 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(G176GAT), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1349GAT) );
  INV_X1 U565 ( .A(n523), .ZN(n584) );
  NAND2_X1 U566 ( .A1(n589), .A2(n584), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n505) );
  XNOR2_X1 U568 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U570 ( .A(G43GAT), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n508), .A2(n587), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(KEYINPUT77), .ZN(n528) );
  AND2_X1 U573 ( .A1(n510), .A2(n528), .ZN(n512) );
  INV_X1 U574 ( .A(KEYINPUT38), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n542) );
  NOR2_X1 U576 ( .A1(n542), .A2(n553), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT40), .B(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1330GAT) );
  AND2_X1 U579 ( .A1(n516), .A2(n295), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT124), .B(n517), .Z(n598) );
  INV_X1 U581 ( .A(n598), .ZN(n594) );
  NAND2_X1 U582 ( .A1(n594), .A2(n587), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n518) );
  XOR2_X1 U584 ( .A(G197GAT), .B(KEYINPUT59), .Z(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1352GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n525) );
  NAND2_X1 U587 ( .A1(n595), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n527) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n546) );
  NAND2_X1 U590 ( .A1(n546), .A2(n528), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n529), .B(KEYINPUT103), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n530), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(KEYINPUT34), .ZN(n532) );
  XNOR2_X1 U594 ( .A(G1GAT), .B(n532), .ZN(G1324GAT) );
  NAND2_X1 U595 ( .A1(n537), .A2(n560), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n535) );
  NAND2_X1 U598 ( .A1(n537), .A2(n562), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G15GAT), .B(n536), .ZN(G1326GAT) );
  NAND2_X1 U601 ( .A1(n564), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U603 ( .A1(n542), .A2(n548), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1328GAT) );
  NOR2_X1 U606 ( .A1(n542), .A2(n551), .ZN(n541) );
  XOR2_X1 U607 ( .A(G36GAT), .B(n541), .Z(G1329GAT) );
  NOR2_X1 U608 ( .A1(n556), .A2(n542), .ZN(n543) );
  XOR2_X1 U609 ( .A(G50GAT), .B(n543), .Z(G1331GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n545) );
  XNOR2_X1 U611 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n548), .A2(n555), .ZN(n549) );
  XOR2_X1 U615 ( .A(n550), .B(n549), .Z(G1332GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n555), .ZN(n552) );
  XOR2_X1 U617 ( .A(G64GAT), .B(n552), .Z(G1333GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n555), .ZN(n554) );
  XOR2_X1 U619 ( .A(G71GAT), .B(n554), .Z(G1334GAT) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n558) );
  XNOR2_X1 U621 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(G78GAT), .B(n559), .ZN(G1335GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n560), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U626 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U628 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n567), .B(n566), .ZN(G1339GAT) );
  NAND2_X1 U631 ( .A1(n587), .A2(n573), .ZN(n569) );
  XOR2_X1 U632 ( .A(G113GAT), .B(KEYINPUT117), .Z(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(G1340GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n571) );
  NAND2_X1 U635 ( .A1(n573), .A2(n423), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G120GAT), .B(n572), .ZN(G1341GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n584), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G134GAT), .B(n576), .ZN(G1343GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n587), .A2(n585), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G141GAT), .B(n579), .ZN(G1344GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n581) );
  NAND2_X1 U646 ( .A1(n585), .A2(n423), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G148GAT), .B(n582), .ZN(G1345GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n595), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U653 ( .A1(n587), .A2(n589), .ZN(n588) );
  XNOR2_X1 U654 ( .A(G169GAT), .B(n588), .ZN(G1348GAT) );
  NAND2_X1 U655 ( .A1(n589), .A2(n595), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U657 ( .A(G204GAT), .B(KEYINPUT61), .Z(n593) );
  NAND2_X1 U658 ( .A1(n591), .A2(n594), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(G1353GAT) );
  XOR2_X1 U660 ( .A(G211GAT), .B(KEYINPUT127), .Z(n597) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n597), .B(n596), .ZN(G1354GAT) );
  NOR2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U664 ( .A(KEYINPUT62), .B(n600), .Z(n601) );
  XNOR2_X1 U665 ( .A(G218GAT), .B(n601), .ZN(G1355GAT) );
endmodule

