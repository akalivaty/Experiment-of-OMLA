//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT68), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT67), .B(G244), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n216), .B(new_n218), .C1(G77), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G87), .A2(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n220), .B(new_n221), .C1(new_n205), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(new_n209), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n203), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n212), .B(new_n225), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT71), .B(KEYINPUT72), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n245), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(new_n227), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n215), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n259), .B(new_n261), .C1(G232), .C2(new_n260), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G97), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT77), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT73), .B(G41), .Z(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI211_X1 g0068(.A(G1), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n255), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n254), .B2(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(G238), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n265), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n275), .B2(new_n277), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n226), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n284), .B1(new_n285), .B2(G68), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n227), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(G68), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT12), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(G13), .A3(G20), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(G68), .ZN(new_n300));
  INV_X1    g0100(.A(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(G68), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(KEYINPUT12), .A3(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n293), .A2(new_n297), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n280), .A2(new_n282), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n278), .A2(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n278), .A2(new_n308), .A3(G169), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n307), .B(new_n309), .C1(new_n310), .C2(new_n278), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n259), .A2(G238), .A3(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n257), .A2(new_n258), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G107), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n270), .ZN(new_n318));
  INV_X1    g0118(.A(new_n269), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n272), .A2(new_n219), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT65), .A2(G20), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT65), .A2(G20), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G77), .ZN(new_n327));
  INV_X1    g0127(.A(new_n283), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n327), .B1(new_n328), .B2(new_n329), .C1(new_n286), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n290), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n294), .A2(G77), .A3(new_n296), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n301), .A2(new_n287), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n269), .B1(new_n317), .B2(new_n270), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n310), .A3(new_n320), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n323), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(KEYINPUT76), .C1(new_n341), .C2(new_n281), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n281), .B1(new_n337), .B2(new_n320), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n336), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(G190), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n312), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n349));
  INV_X1    g0149(.A(G150), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n349), .B1(new_n350), .B2(new_n328), .C1(new_n286), .C2(new_n329), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n290), .B1(new_n214), .B2(new_n301), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n294), .A2(new_n296), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n214), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT9), .ZN(new_n355));
  INV_X1    g0155(.A(G223), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G222), .B2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n255), .B1(new_n259), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n259), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n272), .A2(G226), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n319), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n355), .B(new_n363), .C1(new_n279), .C2(new_n362), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT10), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n362), .A2(G179), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n322), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(new_n354), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n256), .B2(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n257), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n256), .A3(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(G223), .C2(G1698), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n260), .A2(G226), .ZN(new_n377));
  INV_X1    g0177(.A(G87), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n376), .A2(new_n377), .B1(new_n253), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n270), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n272), .A2(G232), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n319), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT81), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(new_n384), .A3(new_n319), .A4(new_n381), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n281), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G190), .B2(new_n382), .ZN(new_n387));
  AND2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(new_n202), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT79), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n375), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n226), .ZN(new_n396));
  AOI21_X1  g0196(.A(G20), .B1(new_n374), .B2(new_n375), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(G68), .C1(new_n397), .C2(new_n395), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT80), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n285), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n302), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT80), .A3(new_n396), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n391), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n294), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n395), .B1(new_n259), .B2(G20), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n315), .A2(new_n226), .A3(KEYINPUT7), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n302), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n391), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n329), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n301), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n353), .B2(new_n412), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n387), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n383), .A2(new_n322), .A3(new_n385), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n382), .A2(G179), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n415), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT18), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n348), .A2(new_n371), .A3(new_n418), .A4(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n294), .B(new_n299), .C1(G1), .C2(new_n253), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G107), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT24), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n374), .A2(G87), .A3(new_n226), .A4(new_n375), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT88), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT22), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n430), .B2(KEYINPUT22), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n315), .A2(new_n326), .A3(KEYINPUT22), .A4(new_n378), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n226), .A2(KEYINPUT23), .A3(G107), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n285), .A2(G33), .A3(G116), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT23), .B1(new_n285), .B2(G107), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n429), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n430), .A2(KEYINPUT22), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT88), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT22), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT24), .B(new_n441), .C1(new_n445), .C2(new_n434), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(new_n290), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n299), .A2(G107), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT25), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G294), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n375), .B1(G250), .B2(G1698), .C1(new_n392), .C2(new_n393), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n260), .A2(G257), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT89), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT89), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n456), .A3(new_n270), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n295), .B(G45), .C1(new_n458), .C2(G41), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT73), .B(G41), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n458), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G274), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n270), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n428), .A2(new_n447), .A3(new_n449), .A4(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n465), .A2(new_n279), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n447), .A2(new_n428), .A3(new_n449), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n322), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n457), .A2(new_n310), .A3(new_n462), .A4(new_n464), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n374), .A2(G68), .A3(new_n226), .A4(new_n375), .ZN(new_n474));
  OAI211_X1 g0274(.A(G33), .B(G97), .C1(new_n324), .C2(new_n325), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(KEYINPUT19), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n324), .B2(new_n325), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n226), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n378), .A2(new_n205), .A3(new_n206), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n290), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n330), .A2(new_n301), .ZN(new_n486));
  INV_X1    g0286(.A(new_n330), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n427), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n295), .A2(G45), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n255), .A2(G250), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G244), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G238), .B2(G1698), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n394), .A2(new_n496), .B1(new_n253), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n493), .B1(new_n498), .B2(new_n270), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n295), .A2(G45), .A3(G274), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(G179), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n270), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n502), .A2(new_n500), .A3(new_n492), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n322), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n485), .A2(new_n505), .A3(new_n486), .A4(new_n488), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n490), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n485), .A2(new_n486), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(G190), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(new_n500), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n427), .A2(G87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n509), .A2(new_n510), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n508), .B1(new_n507), .B2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n427), .A2(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n206), .B1(new_n407), .B2(new_n408), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT6), .B1(new_n207), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n226), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n283), .A2(G77), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT82), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n518), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  OAI221_X1 g0327(.A(new_n517), .B1(G97), .B2(new_n299), .C1(new_n527), .C2(new_n294), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n494), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n260), .A3(new_n257), .A4(new_n258), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n257), .A2(new_n258), .A3(G250), .A4(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n253), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n257), .B2(new_n373), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G244), .A3(new_n260), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(new_n529), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n255), .ZN(new_n539));
  INV_X1    g0339(.A(new_n459), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n267), .B2(KEYINPUT5), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G257), .A3(new_n255), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n462), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n322), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n534), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n394), .A2(new_n494), .A3(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(KEYINPUT4), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n270), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n310), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n528), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n299), .A2(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n407), .A2(new_n408), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G107), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n525), .C1(new_n226), .C2(new_n522), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n554), .B2(new_n290), .ZN(new_n555));
  OAI21_X1  g0355(.A(G200), .B1(new_n539), .B2(new_n543), .ZN(new_n556));
  INV_X1    g0356(.A(new_n543), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(G190), .C1(new_n255), .C2(new_n538), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n555), .A2(new_n517), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n515), .A2(new_n516), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n222), .A2(new_n260), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n536), .B(new_n562), .C1(G264), .C2(new_n260), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n315), .A2(G303), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n255), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n463), .A2(G270), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n322), .B1(new_n567), .B2(new_n462), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n226), .B(new_n532), .C1(G33), .C2(new_n205), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n289), .A2(new_n227), .B1(G20), .B2(new_n497), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT20), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT87), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT87), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n575), .A3(KEYINPUT20), .A4(new_n570), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n426), .A2(KEYINPUT86), .A3(new_n497), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT86), .B1(new_n426), .B2(new_n497), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n301), .A2(new_n497), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT21), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n567), .A2(new_n462), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G200), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n279), .C2(new_n585), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n568), .A2(KEYINPUT21), .A3(new_n582), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n567), .A2(G179), .A3(new_n462), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n584), .A2(new_n588), .A3(new_n589), .A4(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n425), .A2(new_n473), .A3(new_n561), .A4(new_n593), .ZN(G372));
  AND3_X1   g0394(.A1(new_n568), .A2(KEYINPUT21), .A3(new_n582), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n583), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n469), .A2(new_n472), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n560), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n509), .A2(new_n513), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(G200), .B2(new_n511), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n467), .A2(new_n468), .B1(new_n510), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n504), .A2(new_n489), .ZN(new_n603));
  INV_X1    g0403(.A(new_n516), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n605));
  INV_X1    g0405(.A(new_n550), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT26), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n514), .A2(new_n603), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n602), .A2(new_n603), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n425), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n613), .B(KEYINPUT90), .Z(new_n614));
  INV_X1    g0414(.A(new_n370), .ZN(new_n615));
  INV_X1    g0415(.A(new_n424), .ZN(new_n616));
  INV_X1    g0416(.A(new_n305), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n311), .A2(new_n304), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n339), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n616), .B1(new_n621), .B2(new_n418), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n615), .B1(new_n622), .B2(new_n365), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n614), .A2(new_n623), .ZN(G369));
  INV_X1    g0424(.A(G330), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n226), .A2(G13), .ZN(new_n626));
  OR3_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .A3(G1), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT27), .B1(new_n626), .B2(G1), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n593), .B1(new_n587), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n596), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n582), .A3(new_n631), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n625), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n632), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n469), .A2(new_n472), .A3(new_n631), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n467), .A2(new_n468), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n597), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n469), .A2(new_n631), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n637), .B(new_n638), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n473), .A2(new_n634), .A3(new_n632), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n469), .A2(new_n472), .A3(new_n632), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(G399));
  INV_X1    g0447(.A(new_n210), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n460), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G1), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n483), .A2(G116), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n230), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n473), .A2(new_n561), .A3(new_n593), .A4(new_n632), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT30), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n548), .A2(new_n464), .A3(new_n457), .A4(new_n503), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n590), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n457), .A2(new_n503), .A3(new_n464), .ZN(new_n659));
  INV_X1    g0459(.A(new_n462), .ZN(new_n660));
  NOR4_X1   g0460(.A1(new_n565), .A2(new_n566), .A3(new_n310), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(KEYINPUT30), .A3(new_n548), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n548), .A2(new_n503), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n310), .A3(new_n465), .A4(new_n585), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT91), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n631), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(KEYINPUT91), .A3(new_n669), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n655), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT92), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n676), .A3(G330), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n598), .A2(new_n601), .B1(new_n504), .B2(new_n489), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n610), .B1(new_n609), .B2(new_n606), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n515), .A2(new_n516), .A3(new_n550), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n610), .ZN(new_n683));
  AOI211_X1 g0483(.A(new_n679), .B(new_n631), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT29), .B1(new_n612), .B2(new_n632), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n654), .B1(new_n687), .B2(G1), .ZN(G364));
  NOR2_X1   g0488(.A1(G13), .A2(G33), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G20), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n633), .A2(new_n635), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n226), .A2(G190), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n310), .A3(new_n281), .ZN(new_n694));
  INV_X1    g0494(.A(G159), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n279), .A2(new_n281), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n326), .A2(G179), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(G20), .A3(new_n310), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(G50), .B1(G87), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n279), .A2(G179), .A3(G200), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n226), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n205), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n310), .A2(G200), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n693), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n698), .B(new_n707), .C1(G77), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n693), .A2(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n310), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G68), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(G179), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n315), .B1(new_n715), .B2(G107), .ZN(new_n716));
  NOR4_X1   g0516(.A1(new_n226), .A2(new_n310), .A3(new_n279), .A4(G200), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n696), .A2(new_n697), .B1(G58), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n711), .A2(new_n714), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT33), .B(G317), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n713), .A2(new_n720), .B1(G322), .B2(new_n717), .ZN(new_n721));
  INV_X1    g0521(.A(new_n694), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G329), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n315), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n702), .B(KEYINPUT95), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(G303), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n706), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n710), .A2(G311), .B1(G294), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G283), .ZN(new_n730));
  INV_X1    g0530(.A(new_n715), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n727), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G326), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n700), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n719), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n252), .B1(new_n285), .B2(G169), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n231), .A2(new_n268), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n536), .A2(new_n648), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(new_n245), .C2(new_n268), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n259), .A2(G355), .A3(new_n210), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(new_n743), .C1(G116), .C2(new_n210), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n738), .A2(new_n691), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n626), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n651), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n692), .A2(new_n739), .A3(new_n746), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n633), .A2(new_n635), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(G330), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(G396));
  NOR2_X1   g0557(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n612), .A2(new_n632), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n323), .A2(new_n336), .A3(new_n338), .A4(new_n631), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT97), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n631), .A2(new_n336), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n347), .A2(new_n339), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT98), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n762), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n768), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n612), .A2(new_n632), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n678), .A2(KEYINPUT99), .B1(new_n769), .B2(new_n771), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n773), .B(new_n754), .C1(new_n774), .C2(new_n758), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(new_n689), .ZN(new_n776));
  INV_X1    g0576(.A(new_n717), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n731), .A2(new_n378), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(G283), .C2(new_n713), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n726), .A2(G107), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n694), .A2(new_n783), .B1(new_n205), .B2(new_n706), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G303), .B2(new_n701), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n259), .B1(new_n710), .B2(G116), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n781), .A2(new_n782), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n713), .A2(G150), .B1(G143), .B2(new_n717), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n701), .A2(G137), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n695), .C2(new_n709), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT34), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G68), .A2(new_n715), .B1(new_n722), .B2(G132), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n394), .B1(new_n728), .B2(G58), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n725), .A2(new_n214), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n787), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n738), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n738), .A2(new_n689), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT96), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n287), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n776), .A2(new_n750), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n775), .A2(new_n801), .ZN(G384));
  NAND2_X1  g0602(.A1(new_n304), .A2(new_n631), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n312), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n618), .B2(new_n632), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n655), .A2(new_n670), .A3(new_n666), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n770), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n387), .A2(new_n411), .A3(new_n415), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n398), .A2(new_n399), .ZN(new_n811));
  AOI21_X1  g0611(.A(KEYINPUT80), .B1(new_n402), .B2(new_n396), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n390), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n406), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n405), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT100), .B1(new_n815), .B2(new_n415), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT100), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n817), .B(new_n414), .C1(new_n405), .C2(new_n814), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n629), .B1(new_n419), .B2(new_n420), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n810), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT101), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n629), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n422), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n423), .A2(new_n416), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n815), .A2(new_n415), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n817), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n815), .A2(KEYINPUT100), .A3(new_n415), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n820), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n416), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT101), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT37), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n823), .A2(new_n827), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n824), .B(new_n819), .C1(new_n424), .C2(new_n418), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT38), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n809), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT40), .ZN(new_n842));
  INV_X1    g0642(.A(new_n418), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n825), .B1(new_n616), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n826), .B(new_n822), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n840), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n808), .A4(new_n805), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n842), .A2(new_n425), .A3(new_n806), .A4(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(G330), .C1(new_n841), .C2(KEYINPUT40), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n425), .A2(G330), .A3(new_n806), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n619), .A2(new_n632), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n835), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n835), .B2(new_n836), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT39), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n858));
  NAND3_X1  g0658(.A1(new_n846), .A2(new_n840), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n854), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n616), .A2(new_n824), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n339), .A2(new_n631), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n771), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n805), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n839), .B2(new_n840), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n860), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n853), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n425), .A2(new_n686), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n623), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n868), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n295), .B2(new_n747), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT35), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n497), .B1(new_n522), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n229), .B(new_n874), .C1(new_n873), .C2(new_n522), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT36), .ZN(new_n876));
  INV_X1    g0676(.A(G13), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n230), .A2(new_n287), .A3(new_n388), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n201), .A2(new_n302), .ZN(new_n879));
  OAI211_X1 g0679(.A(G1), .B(new_n877), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n876), .A3(new_n880), .ZN(G367));
  NAND4_X1  g0681(.A1(new_n598), .A2(new_n473), .A3(new_n634), .A4(new_n632), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n528), .A2(new_n631), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n550), .A2(new_n559), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n550), .B1(new_n597), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n886), .A2(new_n632), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT43), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n632), .B1(new_n513), .B2(new_n509), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n603), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n609), .B2(new_n889), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT103), .Z(new_n892));
  OAI22_X1  g0692(.A1(new_n883), .A2(new_n887), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n888), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n643), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n606), .A2(new_n631), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n895), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n649), .B(KEYINPUT41), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n642), .A2(new_n644), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n753), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT105), .B1(new_n636), .B2(new_n642), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n905), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n687), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n646), .A2(new_n898), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n646), .A2(new_n898), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT45), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT106), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n686), .ZN(new_n918));
  INV_X1    g0718(.A(new_n677), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n676), .B1(new_n673), .B2(G330), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n909), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n912), .A2(new_n915), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(new_n903), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n902), .B1(new_n926), .B2(new_n687), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n749), .A2(new_n295), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n900), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n754), .B1(new_n892), .B2(new_n691), .ZN(new_n931));
  INV_X1    g0731(.A(new_n741), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n745), .B1(new_n210), .B2(new_n330), .C1(new_n239), .C2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n713), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n695), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n731), .A2(new_n287), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G58), .B2(new_n703), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n259), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n728), .A2(G68), .ZN(new_n940));
  INV_X1    g0740(.A(G143), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n940), .B1(new_n941), .B2(new_n700), .C1(new_n777), .C2(new_n350), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n201), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n939), .B2(new_n942), .C1(new_n944), .C2(new_n709), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT109), .B(G137), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n935), .B(new_n945), .C1(new_n722), .C2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT110), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n715), .A2(G97), .ZN(new_n949));
  INV_X1    g0749(.A(G317), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n394), .C1(new_n950), .C2(new_n694), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT107), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n706), .A2(new_n206), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT46), .B1(new_n703), .B2(G116), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n726), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(G303), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n955), .B1(new_n956), .B2(new_n777), .C1(new_n783), .C2(new_n700), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n730), .B2(new_n709), .C1(new_n778), .C2(new_n934), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n948), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  OAI211_X1 g0761(.A(new_n931), .B(new_n933), .C1(new_n961), .C2(new_n737), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n930), .A2(new_n962), .ZN(G387));
  INV_X1    g0763(.A(new_n922), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n687), .A2(new_n909), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(new_n649), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n909), .A2(new_n929), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT112), .B(G322), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n713), .A2(G311), .B1(new_n701), .B2(new_n968), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n956), .B2(new_n709), .C1(new_n950), .C2(new_n777), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n730), .B2(new_n706), .C1(new_n778), .C2(new_n702), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT49), .Z(new_n973));
  OAI221_X1 g0773(.A(new_n394), .B1(new_n733), .B2(new_n694), .C1(new_n731), .C2(new_n497), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT113), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n949), .B1(new_n214), .B2(new_n777), .C1(new_n695), .C2(new_n700), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n412), .B2(new_n713), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT111), .B(G150), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n722), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n710), .A2(G68), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n728), .A2(new_n487), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n702), .A2(new_n287), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n983), .A2(new_n394), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n738), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n741), .B1(new_n236), .B2(new_n268), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n652), .A2(new_n210), .A3(new_n259), .ZN(new_n988));
  AOI211_X1 g0788(.A(G45), .B(new_n652), .C1(G68), .C2(G77), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n329), .A2(G50), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT50), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n210), .A2(G107), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n745), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n638), .B(new_n691), .C1(new_n640), .C2(new_n641), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n986), .A2(new_n750), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n966), .A2(new_n967), .A3(new_n996), .ZN(G393));
  OAI22_X1  g0797(.A1(new_n777), .A2(new_n783), .B1(new_n950), .B2(new_n700), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT52), .Z(new_n999));
  AOI22_X1  g0799(.A1(new_n722), .A2(new_n968), .B1(G283), .B2(new_n703), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT114), .Z(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(G116), .C2(new_n728), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n778), .B2(new_n709), .C1(new_n956), .C2(new_n934), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n259), .B(new_n1003), .C1(G107), .C2(new_n715), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G159), .A2(new_n717), .B1(new_n701), .B2(G150), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT51), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n394), .B1(new_n710), .B2(new_n412), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n728), .A2(G77), .B1(G68), .B2(new_n703), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n941), .C2(new_n694), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n934), .A2(new_n944), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1006), .A2(new_n1009), .A3(new_n780), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n738), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n250), .A2(new_n741), .B1(G97), .B2(new_n648), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n745), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n750), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n898), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(new_n691), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n924), .A2(new_n896), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n912), .A2(new_n643), .A3(new_n915), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n917), .A2(new_n925), .B1(new_n1022), .B2(new_n964), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1019), .B1(new_n1023), .B2(new_n649), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n928), .B2(new_n1022), .ZN(G390));
  NAND2_X1  g0825(.A1(new_n865), .A2(new_n854), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n857), .A2(new_n859), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT116), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n631), .B(new_n768), .C1(new_n680), .C2(new_n683), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n862), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n680), .A2(new_n683), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n632), .A3(new_n770), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(KEYINPUT116), .A3(new_n863), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1033), .A3(new_n805), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n846), .A2(new_n840), .B1(new_n619), .B2(new_n632), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n678), .A2(new_n770), .A3(new_n805), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1027), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n809), .A2(new_n625), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n929), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n857), .A2(new_n689), .A3(new_n859), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n777), .A2(new_n497), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n713), .A2(G107), .B1(G77), .B2(new_n728), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n730), .B2(new_n700), .C1(new_n778), .C2(new_n694), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G97), .C2(new_n710), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n259), .B1(new_n715), .B2(G68), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n378), .C2(new_n725), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT120), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n703), .A2(new_n979), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT119), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n717), .A2(G132), .ZN(new_n1056));
  INV_X1    g0856(.A(G125), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n694), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n201), .B2(new_n715), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n709), .A2(new_n1061), .B1(new_n695), .B2(new_n706), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n315), .B(new_n1062), .C1(new_n713), .C2(new_n946), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1055), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G128), .B2(new_n701), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n738), .B1(new_n1051), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n799), .A2(new_n329), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1044), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1043), .B1(new_n754), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n623), .A2(new_n851), .A3(new_n869), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n805), .B1(new_n678), .B2(new_n770), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n864), .B1(new_n1071), .B2(new_n1041), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n804), .B1(new_n618), .B2(new_n632), .C1(new_n807), .C2(new_n625), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1037), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1042), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1027), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1041), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT117), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1076), .B(KEYINPUT117), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1077), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1069), .B1(new_n1084), .B2(new_n649), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G378));
  INV_X1    g0886(.A(new_n1070), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT117), .B1(new_n1042), .B2(new_n1076), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1083), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT123), .B1(new_n365), .B2(new_n370), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n354), .A2(new_n824), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n365), .A2(KEYINPUT123), .A3(new_n370), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n842), .A2(G330), .A3(new_n848), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n850), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1102), .A2(new_n867), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n867), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1090), .A2(new_n1107), .A3(KEYINPUT57), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT57), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1070), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1112), .A3(new_n649), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1103), .A2(new_n689), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n984), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n940), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n394), .A2(new_n267), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n713), .A2(G97), .B1(new_n710), .B2(new_n487), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT122), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G116), .C2(new_n701), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n715), .A2(G58), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(KEYINPUT121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1121), .A2(KEYINPUT121), .B1(G283), .B2(new_n722), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1116), .B(new_n1125), .C1(G107), .C2(new_n717), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1117), .B(new_n214), .C1(G33), .C2(G41), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n777), .A2(new_n1130), .B1(new_n350), .B2(new_n706), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n710), .A2(G137), .B1(new_n703), .B2(new_n1060), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1057), .B2(new_n700), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G132), .C2(new_n713), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n722), .A2(G124), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G33), .B(G41), .C1(new_n715), .C2(G159), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n738), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n798), .A2(new_n944), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1114), .A2(new_n750), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1107), .B2(new_n929), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1113), .A2(new_n1144), .ZN(G375));
  NAND2_X1  g0945(.A1(new_n799), .A2(new_n302), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n805), .B2(new_n690), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1123), .B1(new_n934), .B2(new_n1061), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n717), .B2(new_n946), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n694), .A2(new_n1130), .B1(new_n709), .B2(new_n350), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n394), .B(new_n1150), .C1(G132), .C2(new_n701), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n728), .A2(G50), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1121), .A2(KEYINPUT121), .B1(new_n726), .B2(G159), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n982), .B1(new_n956), .B2(new_n694), .C1(new_n934), .C2(new_n497), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n725), .A2(new_n205), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n709), .A2(new_n206), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n777), .A2(new_n730), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n315), .C1(new_n778), .C2(new_n700), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1154), .B1(new_n936), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT124), .Z(new_n1162));
  AOI211_X1 g0962(.A(new_n754), .B(new_n1147), .C1(new_n738), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n929), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1072), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n901), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1167), .B2(new_n1076), .ZN(G381));
  NAND3_X1  g0968(.A1(new_n1113), .A2(new_n1085), .A3(new_n1144), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1169), .A2(G384), .A3(G381), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1022), .A2(new_n928), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n1019), .C1(new_n1023), .C2(new_n649), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n930), .A3(new_n962), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1173), .A2(G396), .A3(G393), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(G407));
  OAI211_X1 g0975(.A(G407), .B(G213), .C1(G343), .C2(new_n1169), .ZN(G409));
  XOR2_X1   g0976(.A(G393), .B(G396), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(G387), .A2(G390), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT127), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n1173), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1179), .B2(new_n1173), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1173), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1172), .B1(new_n962), .B2(new_n930), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT127), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1180), .A3(new_n1173), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1085), .B1(new_n1113), .B2(new_n1144), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1090), .A2(new_n1107), .A3(new_n901), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1085), .A2(new_n1144), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n630), .A2(G213), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT125), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1166), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1164), .A2(new_n1087), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n1070), .A4(new_n1075), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n649), .A4(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(G384), .A3(new_n1165), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G384), .B1(new_n1200), .B2(new_n1165), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1195), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(KEYINPUT125), .A3(new_n1201), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1190), .A2(new_n1194), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1189), .B1(KEYINPUT63), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT63), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT61), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n630), .A2(G213), .A3(G2897), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1205), .B2(new_n1201), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT126), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(KEYINPUT126), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1209), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT62), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n1212), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT61), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1190), .A2(new_n1194), .A3(KEYINPUT62), .A4(new_n1207), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1226), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1189), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1231), .B2(new_n1232), .ZN(G405));
  INV_X1    g1033(.A(new_n1169), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1234), .A2(new_n1190), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1210), .A2(new_n1169), .A3(new_n1212), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(new_n1189), .ZN(G402));
endmodule


