//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT82), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n204), .A2(new_n205), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G148gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n210), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G113gat), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G120gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n231), .A3(new_n229), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n203), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n220), .B(KEYINPUT79), .ZN(new_n237));
  AND2_X1   g036(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n239));
  OAI21_X1  g038(.A(G148gat), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n217), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n206), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n212), .A2(G141gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n207), .B1(new_n217), .B2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n237), .A2(new_n242), .B1(new_n206), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n228), .A2(new_n231), .A3(new_n229), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n231), .B1(new_n228), .B2(new_n229), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT82), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n246), .B2(new_n247), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT80), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n236), .A2(new_n249), .B1(new_n223), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n202), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n223), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n223), .A2(new_n203), .A3(new_n235), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT82), .B1(new_n245), .B2(new_n248), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT83), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n262), .A3(KEYINPUT5), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT84), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n256), .A2(new_n262), .A3(new_n265), .A4(KEYINPUT5), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n258), .B2(new_n259), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n210), .B(new_n269), .C1(new_n218), .C2(new_n222), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n253), .B(new_n270), .C1(new_n271), .C2(new_n245), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n248), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(new_n255), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n264), .A2(new_n266), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n249), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n267), .B1(new_n223), .B2(new_n235), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n276), .A2(new_n272), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(new_n261), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT85), .B(KEYINPUT0), .Z(new_n284));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G57gat), .B(G85gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n290));
  INV_X1    g089(.A(new_n288), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n282), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(KEYINPUT6), .A3(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT75), .B(G8gat), .Z(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT76), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G197gat), .B(G204gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT22), .ZN(new_n303));
  NAND2_X1  g102(.A1(G211gat), .A2(G218gat), .ZN(new_n304));
  OR2_X1    g103(.A1(G211gat), .A2(G218gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT28), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n318), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n320), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n315), .A2(new_n317), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT23), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G169gat), .B2(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT25), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n322), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT67), .A4(new_n333), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n311), .A3(KEYINPUT65), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n325), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n323), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT66), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n342), .A2(new_n344), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n346), .A4(new_n323), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n340), .A2(new_n348), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n336), .A2(KEYINPUT72), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT72), .B1(new_n336), .B2(new_n353), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n310), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT73), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n359), .B(new_n356), .C1(new_n354), .C2(new_n355), .ZN(new_n364));
  INV_X1    g163(.A(new_n310), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n336), .A2(new_n353), .ZN(new_n366));
  INV_X1    g165(.A(new_n356), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n336), .A2(KEYINPUT72), .A3(new_n353), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n360), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n310), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n363), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT74), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n379), .A3(new_n369), .A4(new_n376), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n301), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n374), .B2(new_n310), .ZN(new_n382));
  AOI211_X1 g181(.A(KEYINPUT73), .B(new_n365), .C1(new_n373), .C2(new_n360), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n369), .A4(new_n301), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n363), .A2(new_n369), .A3(new_n376), .A4(new_n301), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n358), .A2(new_n235), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n336), .A2(new_n248), .A3(new_n353), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G227gat), .ZN(new_n394));
  INV_X1    g193(.A(G233gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT64), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT69), .ZN(new_n403));
  INV_X1    g202(.A(G71gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n393), .B2(new_n398), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT34), .B1(new_n393), .B2(new_n396), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n391), .B(new_n392), .C1(new_n394), .C2(new_n395), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n393), .A2(KEYINPUT34), .A3(new_n398), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n410), .B(new_n418), .C1(new_n414), .C2(new_n416), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n408), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n416), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT70), .B1(new_n415), .B2(KEYINPUT34), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n410), .ZN(new_n426));
  INV_X1    g225(.A(new_n408), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n417), .A2(new_n411), .A3(new_n419), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G22gat), .B(G50gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n308), .A2(KEYINPUT88), .A3(new_n302), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n306), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT88), .B1(new_n308), .B2(new_n302), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n359), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n245), .B1(new_n440), .B2(new_n269), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n310), .B1(new_n270), .B2(new_n359), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT89), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(new_n436), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n310), .A2(new_n359), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n245), .B1(new_n448), .B2(new_n271), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n449), .A2(new_n442), .A3(new_n436), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n435), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n434), .B(new_n450), .C1(new_n444), .C2(new_n446), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n431), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n446), .ZN(new_n455));
  INV_X1    g254(.A(new_n269), .ZN(new_n456));
  INV_X1    g255(.A(new_n439), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n306), .A3(new_n437), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n458), .B2(new_n359), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n245), .B2(new_n269), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n459), .A2(new_n245), .B1(new_n460), .B2(new_n310), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n445), .B1(new_n461), .B2(new_n436), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n451), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n434), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n435), .A3(new_n451), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n430), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n422), .A2(new_n429), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n295), .A2(new_n390), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT92), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n295), .A2(new_n468), .A3(new_n390), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n467), .B1(new_n295), .B2(new_n390), .ZN(new_n476));
  INV_X1    g275(.A(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n276), .A2(new_n272), .A3(new_n278), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n261), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT39), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n479), .B(KEYINPUT39), .C1(new_n261), .C2(new_n260), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT40), .A4(new_n291), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n289), .B(new_n482), .C1(new_n381), .C2(new_n389), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n481), .A3(new_n291), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT90), .B(KEYINPUT40), .Z(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT91), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n477), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n293), .A2(new_n294), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n378), .B2(new_n380), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n300), .B1(new_n377), .B2(KEYINPUT37), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n364), .A2(new_n310), .A3(new_n368), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n365), .B2(new_n374), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT38), .B1(new_n496), .B2(KEYINPUT37), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n300), .C1(KEYINPUT37), .C2(new_n377), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n490), .A2(new_n386), .A3(new_n494), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n476), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n501));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n422), .A2(new_n429), .ZN(new_n504));
  MUX2_X1   g303(.A(new_n501), .B(new_n503), .S(new_n504), .Z(new_n505));
  AOI21_X1  g304(.A(new_n475), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(G43gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT15), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT93), .B(G43gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n507), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT15), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n510), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(KEYINPUT16), .A3(new_n525), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(G8gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n529), .A2(G8gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n526), .A2(new_n527), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n535), .A3(new_n521), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n534), .A2(new_n522), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n534), .B(new_n522), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n539), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G113gat), .B(G141gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT11), .B(G169gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n542), .A2(new_n546), .A3(new_n547), .A4(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n559));
  NAND2_X1  g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(KEYINPUT8), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT102), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT96), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(KEYINPUT102), .A3(new_n568), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(KEYINPUT99), .A3(new_n572), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n567), .A2(KEYINPUT99), .A3(new_n568), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n559), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n578), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G230gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(new_n395), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n580), .A2(new_n583), .A3(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n589), .B1(new_n584), .B2(new_n586), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n598), .A2(KEYINPUT103), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT103), .B1(new_n598), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n605));
  NOR2_X1   g404(.A1(new_n578), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n608), .A2(new_n534), .A3(new_n341), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n341), .B1(new_n608), .B2(new_n534), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n534), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G183gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n534), .A3(new_n341), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n614), .A3(new_n606), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT98), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n611), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n611), .B2(new_n615), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G211gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n617), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n615), .A3(new_n618), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n523), .A2(new_n536), .A3(new_n582), .A4(new_n581), .ZN(new_n632));
  AND3_X1   g431(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n522), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n585), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n632), .B2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT100), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n635), .ZN(new_n641));
  INV_X1    g440(.A(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n637), .ZN(new_n645));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(KEYINPUT100), .B(new_n648), .C1(new_n638), .C2(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n652), .A3(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n506), .A2(new_n558), .A3(new_n604), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n490), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  INV_X1    g460(.A(new_n390), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(G8gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n504), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n658), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n505), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n658), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n477), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n476), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n494), .A2(new_n386), .ZN(new_n679));
  INV_X1    g478(.A(new_n498), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n295), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n488), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n467), .B1(new_n682), .B2(new_n483), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n505), .B(new_n678), .C1(new_n681), .C2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n471), .A2(new_n474), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n652), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n604), .A2(new_n558), .ZN(new_n689));
  INV_X1    g488(.A(new_n631), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n517), .A3(new_n490), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n652), .B1(new_n684), .B2(new_n685), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n506), .B2(new_n652), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n691), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(new_n490), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n694), .B1(new_n517), .B2(new_n704), .ZN(G1328gat));
  INV_X1    g504(.A(new_n691), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n699), .A2(new_n518), .A3(new_n662), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n662), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G36gat), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n708), .A2(new_n714), .A3(KEYINPUT46), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n710), .A2(new_n711), .A3(new_n713), .A4(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(new_n511), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n692), .A2(new_n717), .A3(new_n670), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT47), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n703), .B2(new_n672), .ZN(new_n721));
  INV_X1    g520(.A(new_n718), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  NAND2_X1  g524(.A1(new_n703), .A2(new_n477), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n728));
  OR2_X1    g527(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n467), .A2(G50gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n692), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n507), .B1(new_n703), .B2(new_n477), .ZN(new_n734));
  INV_X1    g533(.A(new_n732), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT110), .B(KEYINPUT48), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n733), .A2(new_n736), .ZN(G1331gat));
  NOR4_X1   g536(.A1(new_n506), .A2(new_n557), .A3(new_n603), .A4(new_n657), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n490), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT111), .B(G57gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n662), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  NAND2_X1  g544(.A1(new_n738), .A2(new_n670), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n404), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n738), .A2(G71gat), .A3(new_n672), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n738), .A2(new_n477), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n631), .A2(new_n557), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n603), .B(new_n754), .C1(new_n701), .C2(new_n702), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(G85gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n686), .A2(new_n687), .A3(new_n753), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n490), .A3(new_n604), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n756), .A2(new_n490), .B1(new_n561), .B2(new_n762), .ZN(G1336gat));
  NAND2_X1  g562(.A1(new_n701), .A2(new_n702), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(new_n604), .A3(new_n662), .A4(new_n753), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n761), .A2(new_n562), .A3(new_n604), .A4(new_n662), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1337gat));
  AND2_X1   g571(.A1(new_n755), .A2(new_n672), .ZN(new_n773));
  INV_X1    g572(.A(new_n761), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n504), .A2(G99gat), .A3(new_n603), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT112), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n773), .A2(new_n406), .B1(new_n774), .B2(new_n776), .ZN(G1338gat));
  NOR2_X1   g576(.A1(new_n467), .A2(G106gat), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n506), .A2(new_n758), .A3(new_n652), .A4(new_n754), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n699), .B2(new_n753), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n604), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n761), .A2(KEYINPUT113), .A3(new_n604), .A4(new_n778), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n755), .B2(new_n477), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n764), .A2(new_n604), .A3(new_n753), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n789), .B2(new_n467), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n761), .A2(new_n793), .A3(new_n604), .A4(new_n778), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n795), .ZN(G1339gat));
  NAND2_X1  g595(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT118), .B(G113gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n601), .A2(new_n557), .A3(new_n602), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n655), .A2(new_n656), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n543), .A2(new_n545), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n552), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n556), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n601), .B2(new_n602), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n584), .A2(new_n589), .A3(new_n586), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n591), .A2(new_n807), .A3(KEYINPUT54), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n599), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n596), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n557), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n598), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n806), .B(new_n652), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n805), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n687), .B1(new_n817), .B2(new_n815), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n690), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n655), .A2(new_n820), .A3(new_n799), .A4(new_n656), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AND4_X1   g621(.A1(new_n490), .A2(new_n822), .A3(new_n390), .A4(new_n468), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n557), .ZN(new_n824));
  MUX2_X1   g623(.A(new_n797), .B(new_n798), .S(new_n824), .Z(G1340gat));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n604), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n631), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n687), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(G134gat), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT56), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(G134gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1343gat));
  NAND3_X1  g633(.A1(new_n505), .A2(new_n490), .A3(new_n390), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n822), .A2(new_n477), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n477), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n835), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n477), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n822), .B2(new_n477), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n841), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n557), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n238), .A2(new_n239), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n558), .B1(new_n853), .B2(new_n846), .ZN(new_n854));
  INV_X1    g653(.A(new_n850), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT120), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n836), .A2(new_n835), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n216), .A3(new_n557), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n851), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n850), .B1(new_n852), .B2(new_n558), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(G1344gat));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n842), .A2(new_n847), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n603), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n819), .A2(new_n800), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n837), .B1(new_n868), .B2(new_n467), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n603), .B1(new_n869), .B2(new_n839), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(KEYINPUT59), .A3(new_n843), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n212), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G148gat), .B1(new_n857), .B2(new_n604), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(KEYINPUT59), .B2(new_n873), .ZN(G1345gat));
  AOI21_X1  g673(.A(G155gat), .B1(new_n857), .B2(new_n631), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n866), .A2(new_n690), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n857), .B2(new_n687), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n866), .A2(new_n652), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(G162gat), .ZN(G1347gat));
  NAND2_X1  g679(.A1(new_n662), .A2(new_n295), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n504), .A3(new_n477), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n822), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n558), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n328), .ZN(G1348gat));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n603), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(new_n329), .ZN(G1349gat));
  INV_X1    g686(.A(new_n883), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n631), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G183gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n312), .A2(new_n313), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n889), .ZN(new_n892));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1350gat));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n687), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(G190gat), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(G190gat), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT61), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n836), .A2(new_n672), .A3(new_n881), .ZN(new_n901));
  XOR2_X1   g700(.A(KEYINPUT123), .B(G197gat), .Z(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n557), .A3(new_n902), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n672), .B(new_n881), .C1(new_n869), .C2(new_n839), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n557), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT124), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n902), .ZN(G1352gat));
  INV_X1    g706(.A(new_n901), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(G204gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n603), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT126), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n870), .A2(new_n295), .A3(new_n505), .A4(new_n662), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n909), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(G1353gat));
  NAND2_X1  g715(.A1(new_n904), .A2(new_n631), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G211gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT63), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n908), .A2(G211gat), .A3(new_n690), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(G1354gat));
  INV_X1    g720(.A(G218gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n922), .A3(new_n687), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n904), .A2(new_n687), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(G1355gat));
endmodule


