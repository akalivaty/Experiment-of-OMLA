//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G107), .C2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n204), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n225), .A2(new_n210), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n209), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G222), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n256), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n262), .C1(G77), .C2(new_n255), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n260), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(new_n203), .C1(G41), .C2(G45), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n261), .A2(new_n267), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n263), .B(new_n271), .C1(new_n221), .C2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(G179), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n230), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G50), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n281), .A2(new_n204), .A3(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n220), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(KEYINPUT8), .A2(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT8), .A2(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n204), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n288), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n277), .A2(new_n230), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n280), .B(new_n283), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n273), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n274), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n273), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n300), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n273), .A2(G200), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n307), .A3(new_n311), .ZN(new_n313));
  INV_X1    g0113(.A(new_n310), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT10), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n303), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT16), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n255), .B2(G20), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n210), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G58), .A2(G68), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n233), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n286), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n317), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT7), .B1(new_n322), .B2(new_n204), .ZN(new_n334));
  NOR4_X1   g0134(.A1(new_n320), .A2(new_n321), .A3(new_n318), .A4(G20), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n329), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT16), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n338), .A3(new_n278), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n281), .A2(G1), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n292), .A2(new_n342), .A3(new_n294), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n279), .B1(new_n292), .B2(new_n294), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n292), .A2(new_n294), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT74), .B(new_n343), .C1(new_n347), .C2(new_n279), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n258), .A2(new_n256), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n221), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(new_n320), .C2(new_n321), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n262), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n272), .A2(new_n226), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n357), .A3(new_n271), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G200), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n261), .B1(new_n352), .B2(new_n353), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n360), .A2(new_n361), .A3(new_n356), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G190), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n339), .A2(new_n349), .A3(new_n359), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n339), .A2(new_n349), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n355), .A2(new_n357), .A3(new_n368), .A4(new_n271), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n362), .B2(G169), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT18), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT18), .B1(new_n367), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT75), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n367), .A2(new_n371), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT18), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n366), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n299), .B2(new_n342), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n282), .A2(new_n278), .A3(KEYINPUT68), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n276), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G20), .A2(G77), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n388), .B2(new_n296), .C1(new_n287), .C2(new_n291), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n386), .A2(G77), .B1(new_n278), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n282), .A2(new_n222), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT69), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT69), .A3(new_n391), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G238), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n255), .B(new_n394), .C1(new_n226), .C2(G1698), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n395), .B(new_n262), .C1(G107), .C2(new_n255), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n271), .C1(new_n223), .C2(new_n272), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G200), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n393), .B(new_n398), .C1(new_n306), .C2(new_n397), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n316), .B(new_n381), .C1(new_n392), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n221), .A2(new_n256), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(G232), .B2(new_n256), .C1(new_n320), .C2(new_n321), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n361), .B1(new_n262), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n261), .A2(G238), .A3(new_n267), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT3), .ZN(new_n409));
  INV_X1    g0209(.A(G33), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT3), .A2(G33), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(new_n412), .B1(new_n226), .B2(G1698), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n402), .B1(G33), .B2(G97), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n271), .B(new_n407), .C1(new_n414), .C2(new_n261), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(G169), .C1(new_n408), .C2(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n406), .A2(new_n401), .A3(new_n407), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G179), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT72), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .A4(G179), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n418), .A2(new_n420), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n282), .A2(KEYINPUT70), .A3(new_n210), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT12), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT70), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n342), .B2(G68), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n429), .B(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n222), .B2(new_n296), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n434), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT11), .B1(new_n434), .B2(new_n278), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G68), .B(new_n275), .C1(new_n383), .C2(new_n384), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n427), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  INV_X1    g0241(.A(new_n439), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n421), .A2(new_n422), .A3(G190), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n421), .B2(new_n422), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(KEYINPUT71), .A3(new_n442), .A4(new_n443), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n390), .A2(new_n391), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n397), .A2(G179), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n397), .A2(new_n301), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n440), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n261), .A2(G274), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G41), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(G41), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(KEYINPUT78), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n458), .A2(new_n459), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n261), .A2(new_n462), .A3(G274), .A4(new_n457), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n461), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n460), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT79), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n215), .A2(G1698), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n474), .B1(G250), .B2(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n410), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n262), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n457), .A2(new_n470), .A3(new_n469), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G264), .A3(new_n261), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT86), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(new_n482), .A3(G264), .A4(new_n261), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n473), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G179), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n473), .A2(new_n480), .A3(new_n478), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G169), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT83), .A2(G87), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n204), .B(new_n495), .C1(new_n320), .C2(new_n321), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT22), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n255), .A2(new_n498), .A3(new_n204), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n410), .A2(new_n249), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n204), .A2(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT23), .ZN(new_n506));
  AND4_X1   g0306(.A1(new_n494), .A2(new_n500), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n503), .B1(new_n497), .B2(new_n499), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n494), .B1(new_n508), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n493), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n278), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n341), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n203), .A2(G33), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n299), .A2(new_n342), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n247), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n490), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n517), .ZN(new_n519));
  AOI211_X1 g0319(.A(KEYINPUT85), .B(new_n519), .C1(new_n510), .C2(new_n278), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n489), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n500), .A2(new_n504), .A3(new_n506), .ZN(new_n522));
  INV_X1    g0322(.A(new_n494), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n508), .A2(new_n494), .A3(new_n506), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n492), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n517), .B1(new_n526), .B2(new_n299), .ZN(new_n527));
  INV_X1    g0327(.A(new_n487), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n473), .A2(new_n484), .A3(new_n478), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n306), .B1(new_n529), .B2(new_n445), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n256), .C1(new_n320), .C2(new_n321), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n533), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n255), .A2(G244), .A3(new_n256), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n262), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n479), .A2(new_n261), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G257), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n473), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n515), .A2(new_n214), .ZN(new_n545));
  OAI21_X1  g0345(.A(G107), .B1(new_n334), .B2(new_n335), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n286), .A2(G77), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n214), .A2(new_n247), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n546), .B(new_n547), .C1(new_n204), .C2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n545), .B1(new_n554), .B2(new_n278), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n342), .A2(G97), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT76), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n540), .A2(new_n473), .A3(G190), .A4(new_n542), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n544), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n545), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n247), .B1(new_n319), .B2(new_n323), .ZN(new_n561));
  INV_X1    g0361(.A(new_n547), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n204), .B1(new_n551), .B2(new_n552), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n560), .B(new_n557), .C1(new_n564), .C2(new_n299), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n543), .A2(new_n301), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n540), .A2(new_n473), .A3(new_n368), .A4(new_n542), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n531), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n541), .A2(G270), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n256), .A2(G257), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G264), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n320), .C2(new_n321), .ZN(new_n574));
  INV_X1    g0374(.A(G303), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n411), .A2(new_n575), .A3(new_n412), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n262), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n473), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G116), .B(new_n514), .C1(new_n383), .C2(new_n384), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n341), .A2(G20), .A3(new_n249), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n537), .B(new_n204), .C1(G33), .C2(new_n214), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n249), .A2(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n278), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n278), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n578), .A2(new_n588), .A3(G169), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT21), .ZN(new_n590));
  INV_X1    g0390(.A(new_n577), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n467), .B2(new_n472), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n592), .A2(G179), .A3(new_n571), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n589), .A2(new_n590), .B1(new_n593), .B2(new_n588), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n578), .A2(new_n588), .A3(KEYINPUT21), .A4(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n301), .B1(new_n592), .B2(new_n571), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n588), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n578), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n588), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n306), .C2(new_n578), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n594), .A2(new_n597), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n204), .B1(new_n404), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G87), .ZN(new_n606));
  AND4_X1   g0406(.A1(KEYINPUT80), .A2(new_n606), .A3(new_n214), .A4(new_n247), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G87), .A2(G97), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT80), .B1(new_n608), .B2(new_n247), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n604), .B1(new_n296), .B2(new_n214), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n255), .A2(new_n204), .A3(G68), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n278), .ZN(new_n614));
  INV_X1    g0414(.A(new_n515), .ZN(new_n615));
  INV_X1    g0415(.A(new_n388), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n388), .A2(new_n282), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n211), .A2(new_n256), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n223), .A2(G1698), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n320), .C2(new_n321), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n261), .B1(new_n622), .B2(new_n502), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n261), .B(G250), .C1(G1), .C2(new_n456), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n623), .A2(new_n625), .A3(new_n458), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n368), .ZN(new_n627));
  INV_X1    g0427(.A(new_n458), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n411), .A2(new_n412), .B1(new_n223), .B2(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n501), .B1(new_n629), .B2(new_n620), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n624), .C1(new_n630), .C2(new_n261), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n301), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n619), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(G190), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(G200), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n613), .A2(new_n278), .B1(new_n282), .B2(new_n388), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n615), .A2(G87), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT81), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n633), .B2(new_n638), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n521), .A2(new_n570), .A3(new_n603), .A4(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n400), .A2(new_n455), .A3(new_n643), .ZN(G372));
  AOI21_X1  g0444(.A(new_n454), .B1(new_n447), .B2(new_n449), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n440), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n427), .A2(new_n439), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT89), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  INV_X1    g0450(.A(new_n366), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n377), .A2(new_n379), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n312), .A2(new_n315), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n303), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n400), .A2(new_n455), .ZN(new_n657));
  INV_X1    g0457(.A(new_n633), .ZN(new_n658));
  INV_X1    g0458(.A(new_n634), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(KEYINPUT87), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n635), .A2(new_n636), .A3(new_n662), .A4(new_n637), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(new_n568), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n633), .B(KEYINPUT88), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n640), .A2(new_n641), .A3(new_n568), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n665), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n485), .A2(G200), .B1(G190), .B2(new_n487), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n511), .A2(new_n671), .A3(new_n517), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n664), .A2(new_n672), .A3(new_n568), .A4(new_n559), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n589), .A2(new_n590), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n593), .A2(new_n588), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n597), .A2(new_n674), .A3(new_n599), .A4(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n511), .A2(new_n517), .B1(new_n488), .B2(new_n486), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n657), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n656), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n521), .A2(new_n672), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n527), .A2(KEYINPUT85), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n511), .A2(new_n490), .A3(new_n517), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n341), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .A3(G20), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT27), .B1(new_n687), .B2(G20), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n683), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n692), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n521), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n603), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n601), .A2(new_n694), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n676), .B2(new_n698), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n701), .A3(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n677), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n678), .B1(new_n683), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n694), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n207), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OR3_X1    g0509(.A1(new_n607), .A2(new_n609), .A3(G116), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n234), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(new_n668), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n664), .A2(new_n666), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT26), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n669), .A2(new_n665), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n676), .B1(new_n686), .B2(new_n489), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n673), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n715), .B1(new_n721), .B2(new_n694), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n715), .B(new_n694), .C1(new_n670), .C2(new_n679), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n540), .A2(new_n473), .A3(new_n542), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n593), .A2(new_n726), .A3(new_n485), .A4(new_n626), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n543), .A2(new_n368), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n529), .A3(new_n578), .A4(new_n631), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n578), .A2(new_n368), .A3(new_n631), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n485), .A4(new_n726), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n692), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n737), .A3(new_n692), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n633), .A2(new_n638), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT81), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n531), .A3(new_n569), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n521), .A3(new_n603), .A4(new_n694), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n725), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n722), .A2(new_n724), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n714), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n281), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n709), .A2(G1), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT90), .Z(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n701), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n230), .B1(G20), .B2(new_n301), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n253), .A2(G45), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n707), .A2(new_n255), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n761), .B(new_n762), .C1(G45), .C2(new_n234), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n207), .A2(new_n255), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n763), .B1(G116), .B2(new_n207), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n753), .B(new_n758), .C1(new_n760), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n204), .A2(new_n368), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n445), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n204), .A2(G179), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n779), .A2(new_n776), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(G329), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT93), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  INV_X1    g0586(.A(new_n769), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n306), .A3(new_n445), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n781), .B1(new_n575), .B2(new_n785), .C1(new_n786), .C2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n787), .A2(new_n306), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(new_n770), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n306), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n204), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n322), .B1(new_n799), .B2(new_n476), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n790), .A2(new_n794), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n777), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n791), .A2(G58), .B1(G77), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT92), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n804), .B(new_n255), .C1(new_n220), .C2(new_n789), .ZN(new_n805));
  INV_X1    g0605(.A(new_n795), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G68), .A2(new_n772), .B1(new_n806), .B2(G107), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n807), .B1(new_n214), .B2(new_n799), .C1(new_n785), .C2(new_n606), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n780), .A2(G159), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n805), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n759), .B1(new_n801), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n700), .A2(new_n725), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n752), .B1(new_n701), .B2(G330), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n768), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n680), .A2(new_n694), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n451), .A2(new_n692), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT95), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT95), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n451), .A2(new_n820), .A3(new_n692), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(new_n399), .C2(new_n392), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n454), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n454), .A2(new_n692), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n824), .B1(new_n822), .B2(new_n454), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n694), .B(new_n828), .C1(new_n670), .C2(new_n679), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(new_n746), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n753), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n795), .A2(new_n210), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n791), .A2(G143), .B1(G150), .B2(new_n772), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G159), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n789), .C1(new_n836), .C2(new_n777), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  INV_X1    g0639(.A(new_n799), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n833), .B(new_n839), .C1(G58), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n785), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G50), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n322), .B1(new_n838), .B2(KEYINPUT34), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G132), .B2(new_n780), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n789), .A2(new_n575), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n840), .A2(G97), .B1(new_n772), .B2(G283), .ZN(new_n848));
  INV_X1    g0648(.A(new_n780), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n775), .B2(new_n849), .C1(new_n476), .C2(new_n792), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n847), .B(new_n850), .C1(G116), .C2(new_n802), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n255), .B1(new_n806), .B2(G87), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n247), .C2(new_n785), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT94), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n759), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n826), .A2(new_n754), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n759), .A2(new_n754), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n222), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n752), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  AND3_X1   g0660(.A1(new_n734), .A2(new_n737), .A3(new_n692), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n737), .B1(new_n734), .B2(new_n692), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n643), .A2(new_n692), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n739), .A2(new_n745), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n364), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n339), .A2(new_n349), .B1(new_n370), .B2(new_n690), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n690), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n367), .B1(new_n371), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n364), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT96), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n870), .B2(new_n874), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n367), .A2(new_n871), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(KEYINPUT38), .C1(new_n381), .C2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n374), .A2(new_n380), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n882), .B2(new_n651), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(new_n872), .B2(new_n364), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT96), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n439), .A2(new_n692), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n440), .A2(new_n450), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n440), .A2(new_n450), .ZN(new_n893));
  INV_X1    g0693(.A(new_n891), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n826), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n867), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n879), .B1(new_n651), .B2(new_n653), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n884), .A2(new_n885), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n881), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n880), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n867), .A2(KEYINPUT40), .A3(new_n903), .A4(new_n896), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n867), .A2(new_n657), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n905), .B(new_n906), .Z(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n440), .A2(new_n450), .A3(new_n891), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n891), .B1(new_n440), .B2(new_n450), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n829), .B2(new_n825), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n890), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n653), .A2(new_n871), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT97), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT97), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n913), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n440), .A2(new_n692), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n887), .B(new_n886), .C1(new_n381), .C2(new_n879), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n902), .B(new_n922), .C1(new_n923), .C2(new_n881), .ZN(new_n924));
  AOI22_X1  g0724(.A1(KEYINPUT98), .A2(new_n924), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n890), .A2(KEYINPUT98), .A3(KEYINPUT39), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n921), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n908), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n657), .B1(new_n722), .B2(new_n724), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n656), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n930), .B(new_n932), .Z(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n203), .B2(new_n749), .ZN(new_n934));
  INV_X1    g0734(.A(new_n553), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n249), .B1(new_n935), .B2(KEYINPUT35), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n232), .C1(KEYINPUT35), .C2(new_n935), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  AND4_X1   g0738(.A1(G77), .A2(new_n235), .A3(new_n327), .A4(new_n328), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n210), .A2(G50), .ZN(new_n940));
  OAI211_X1 g0740(.A(G1), .B(new_n281), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n676), .A2(new_n694), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n693), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n694), .B1(new_n555), .B2(new_n557), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n569), .A2(KEYINPUT100), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT100), .B1(new_n569), .B2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n945), .A2(KEYINPUT42), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n568), .B1(new_n950), .B2(new_n521), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n694), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT42), .B1(new_n945), .B2(new_n950), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n694), .B1(new_n636), .B2(new_n637), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n664), .B(new_n716), .S(new_n956), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n693), .A2(new_n695), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n960), .A2(new_n700), .A3(new_n725), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n950), .B1(new_n568), .B2(new_n694), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n955), .A2(new_n963), .A3(new_n958), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n708), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n960), .B1(new_n700), .B2(new_n725), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n702), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n944), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n704), .A2(new_n950), .A3(new_n694), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n962), .A2(new_n705), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n961), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n978), .B(KEYINPUT45), .Z(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n976), .A3(new_n702), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n974), .A2(new_n980), .A3(new_n982), .A4(new_n747), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n971), .B1(new_n983), .B2(new_n747), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n750), .A2(G1), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n969), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n785), .A2(new_n225), .B1(new_n835), .B2(new_n849), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT102), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n840), .A2(G68), .B1(new_n772), .B2(G159), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n220), .B2(new_n777), .ZN(new_n990));
  INV_X1    g0790(.A(G143), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n789), .A2(new_n991), .B1(new_n795), .B2(new_n222), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n990), .A2(new_n992), .A3(new_n322), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n988), .B(new_n993), .C1(new_n285), .C2(new_n792), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n795), .A2(new_n214), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n792), .A2(new_n575), .B1(new_n247), .B2(new_n799), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(G311), .C2(new_n788), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n842), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT101), .B(G317), .Z(new_n999));
  AOI21_X1  g0799(.A(new_n255), .B1(new_n780), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n796), .B2(new_n777), .C1(new_n476), .C2(new_n771), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT46), .B1(new_n842), .B2(G116), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n759), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n957), .A2(new_n757), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n762), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n760), .B1(new_n207), .B2(new_n388), .C1(new_n239), .C2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n752), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n986), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT103), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT103), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n986), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(G387));
  OR2_X1    g0815(.A1(new_n974), .A2(new_n747), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n974), .A2(new_n747), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n708), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n974), .A2(new_n985), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n840), .A2(new_n616), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n285), .B2(new_n849), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n322), .B(new_n1021), .C1(G50), .C2(new_n791), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n802), .A2(G68), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n295), .A2(new_n772), .B1(new_n788), .B2(G159), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n995), .B1(new_n842), .B2(G77), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n788), .A2(G322), .B1(G311), .B2(new_n772), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT106), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n791), .A2(new_n999), .B1(G303), .B2(new_n802), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n796), .B2(new_n799), .C1(new_n476), .C2(new_n785), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT49), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n322), .B1(new_n249), .B2(new_n795), .C1(new_n849), .C2(new_n786), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1026), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1035), .A2(new_n759), .B1(new_n960), .B2(new_n756), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n762), .B1(new_n244), .B2(new_n456), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n711), .B2(new_n766), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n291), .A2(G50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n711), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1038), .A2(new_n1043), .B1(new_n247), .B2(new_n707), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n760), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n752), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT105), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n1036), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1018), .A2(new_n1019), .A3(new_n1048), .ZN(G393));
  NAND2_X1  g0849(.A1(new_n980), .A2(new_n982), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1017), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(new_n708), .A3(new_n983), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n980), .A2(new_n982), .A3(new_n985), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n760), .B1(new_n214), .B2(new_n207), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n250), .B2(new_n762), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n791), .A2(G159), .B1(new_n788), .B2(G150), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT51), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n255), .B1(new_n777), .B2(new_n291), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G77), .B2(new_n840), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n849), .A2(new_n991), .B1(new_n606), .B2(new_n795), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G50), .B2(new_n772), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n842), .A2(G68), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT107), .Z(new_n1064));
  OAI21_X1  g0864(.A(new_n322), .B1(new_n849), .B2(new_n793), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n791), .A2(G311), .B1(new_n788), .B2(G317), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(G107), .C2(new_n806), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n796), .B2(new_n785), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G294), .A2(new_n802), .B1(new_n772), .B2(G303), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n249), .B2(new_n799), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT108), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n753), .B(new_n1055), .C1(new_n1073), .C2(new_n759), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n962), .B2(new_n757), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1052), .A2(new_n1053), .A3(new_n1075), .ZN(G390));
  NAND4_X1  g0876(.A1(new_n864), .A2(G330), .A3(new_n866), .A4(new_n828), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n911), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n721), .A2(new_n694), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n824), .B1(new_n1079), .B2(new_n823), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n895), .A2(new_n892), .ZN(new_n1081));
  AND4_X1   g0881(.A1(G330), .A2(new_n863), .A3(new_n1081), .A4(new_n828), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n864), .A2(new_n896), .A3(new_n866), .A4(G330), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n863), .A2(G330), .A3(new_n828), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n911), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n829), .A2(new_n825), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n864), .A2(new_n657), .A3(new_n866), .A4(G330), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n656), .A2(new_n931), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT109), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT109), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1096), .B(new_n1093), .C1(new_n1084), .C2(new_n1090), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n924), .A2(KEYINPUT98), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n882), .A2(new_n651), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n879), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT38), .B1(new_n1102), .B2(new_n878), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n883), .A2(new_n888), .A3(new_n881), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT39), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1099), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1089), .A2(new_n1081), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n921), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n926), .A3(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n903), .C1(new_n1080), .C2(new_n911), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1085), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1083), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT110), .B1(new_n1098), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1082), .B1(new_n1077), .B2(new_n911), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n1080), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n1093), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1110), .A2(new_n1082), .A3(new_n1111), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1085), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1096), .B1(new_n1117), .B2(new_n1093), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1091), .A2(KEYINPUT109), .A3(new_n1094), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT110), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1115), .A2(new_n708), .A3(new_n1122), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1106), .A2(new_n754), .A3(new_n926), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n759), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n322), .B1(new_n222), .B2(new_n799), .C1(new_n785), .C2(new_n606), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n833), .B(new_n1132), .C1(G116), .C2(new_n791), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n788), .A2(G283), .B1(G97), .B2(new_n802), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n247), .B2(new_n771), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT112), .Z(new_n1136));
  OAI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(new_n476), .C2(new_n849), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n322), .B1(new_n780), .B2(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n220), .B2(new_n795), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT111), .Z(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G132), .B2(new_n791), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n802), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n788), .A2(G128), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n799), .A2(new_n836), .B1(new_n771), .B2(new_n835), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n842), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT53), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n785), .B2(new_n285), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1131), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n753), .B(new_n1151), .C1(new_n347), .C2(new_n857), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1114), .A2(new_n985), .B1(new_n1130), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1129), .A2(new_n1153), .ZN(G378));
  NAND2_X1  g0954(.A1(new_n1122), .A2(new_n1094), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n300), .A2(new_n871), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n316), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n316), .A2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT117), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n918), .B1(new_n913), .B2(new_n915), .ZN(new_n1168));
  AOI211_X1 g0968(.A(KEYINPUT97), .B(new_n914), .C1(new_n912), .C2(new_n890), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1108), .B1(new_n1106), .B2(new_n926), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1167), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n920), .A2(new_n928), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n899), .A2(G330), .A3(new_n904), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1155), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n708), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n799), .A2(new_n210), .B1(new_n777), .B2(new_n388), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G41), .B(new_n255), .C1(new_n780), .C2(G283), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n225), .B2(new_n795), .C1(new_n785), .C2(new_n222), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT113), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(G116), .C2(new_n788), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n214), .B2(new_n771), .C1(new_n247), .C2(new_n792), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT58), .Z(new_n1187));
  NAND2_X1  g0987(.A1(new_n842), .A2(new_n1142), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n772), .A2(G132), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n791), .A2(G128), .B1(G137), .B2(new_n802), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G125), .A2(new_n788), .B1(new_n840), .B2(G150), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n410), .B(new_n463), .C1(new_n795), .C2(new_n836), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G124), .B2(new_n780), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n220), .B1(new_n320), .B2(G41), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n759), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n857), .A2(new_n220), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n752), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n755), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1170), .A2(new_n1171), .A3(new_n1167), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1173), .B1(new_n920), .B2(new_n928), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1175), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(KEYINPUT118), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1122), .B2(new_n1094), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n985), .B1(new_n1214), .B2(new_n708), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1180), .B(new_n1205), .C1(new_n1213), .C2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1117), .A2(new_n1093), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1125), .A2(new_n970), .A3(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n785), .A2(new_n214), .B1(new_n575), .B2(new_n849), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT121), .Z(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1020), .C1(new_n796), .C2(new_n792), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n788), .A2(G294), .B1(G107), .B2(new_n802), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n249), .B2(new_n771), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT119), .Z(new_n1224));
  OAI21_X1  g1024(.A(new_n322), .B1(new_n795), .B2(new_n222), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT120), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1221), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT122), .Z(new_n1228));
  NOR2_X1   g1028(.A1(new_n785), .A2(new_n836), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n795), .A2(new_n225), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n322), .B1(new_n780), .B2(G128), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n285), .B2(new_n777), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G137), .C2(new_n791), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n788), .A2(G132), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n840), .A2(G50), .B1(new_n772), .B2(new_n1142), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n753), .B1(new_n1237), .B2(new_n759), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n755), .B2(new_n1081), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n210), .B2(new_n857), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1091), .B2(new_n985), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1218), .A2(new_n1241), .ZN(G381));
  NOR3_X1   g1042(.A1(new_n1177), .A2(new_n1178), .A3(new_n1206), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT118), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1214), .A2(new_n708), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n985), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1204), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1129), .A2(new_n1153), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1180), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1251), .A2(G390), .A3(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1251), .ZN(G409));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G343), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G2897), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n832), .A2(new_n859), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1084), .A2(new_n1090), .A3(KEYINPUT60), .A4(new_n1093), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT123), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1117), .A2(new_n1264), .A3(KEYINPUT60), .A4(new_n1093), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n709), .B1(new_n1217), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1118), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(KEYINPUT124), .B(new_n1261), .C1(new_n1270), .C2(new_n1241), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G384), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1261), .A2(KEYINPUT124), .ZN(new_n1274));
  AND4_X1   g1074(.A1(new_n1241), .A2(new_n1270), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1260), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1270), .A2(new_n1241), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1272), .A3(G384), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1270), .A2(new_n1274), .A3(new_n1241), .A4(new_n1273), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(G2897), .A3(new_n1279), .A4(new_n1259), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1204), .B1(new_n1282), .B2(new_n985), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1129), .A2(new_n1283), .A3(new_n1153), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1207), .A2(new_n1212), .A3(new_n970), .A4(new_n1155), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1259), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G375), .A2(G378), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1257), .B1(new_n1288), .B2(KEYINPUT61), .ZN(new_n1289));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n986), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1013), .B1(new_n986), .B2(new_n1010), .ZN(new_n1292));
  OAI211_X1 g1092(.A(KEYINPUT126), .B(new_n1290), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1252), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G390), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n986), .A2(G390), .A3(new_n1010), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT126), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1293), .B(new_n1295), .C1(new_n1296), .C2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1011), .A2(new_n1290), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1297), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1252), .A3(new_n1294), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1250), .B1(new_n1249), .B2(new_n1180), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1285), .A2(new_n1129), .A3(new_n1153), .A4(new_n1283), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1259), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1304), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(KEYINPUT127), .A3(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1289), .A2(new_n1303), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1287), .A2(new_n1313), .A3(new_n1307), .A4(new_n1306), .ZN(new_n1314));
  XOR2_X1   g1114(.A(new_n1314), .B(KEYINPUT62), .Z(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1286), .A2(new_n1317), .A3(new_n1313), .A4(new_n1287), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT125), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT125), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1286), .A2(new_n1321), .A3(new_n1287), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1304), .A3(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(new_n1310), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1312), .A2(new_n1315), .B1(new_n1324), .B2(new_n1325), .ZN(G405));
  AOI21_X1  g1126(.A(new_n1313), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1299), .A2(new_n1302), .A3(new_n1313), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1328), .A2(new_n1329), .B1(new_n1251), .B2(new_n1287), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1329), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1251), .A2(new_n1287), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1331), .A2(new_n1327), .A3(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1330), .A2(new_n1333), .ZN(G402));
endmodule


