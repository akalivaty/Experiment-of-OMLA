

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U556 ( .A(n958), .ZN(n781) );
  XNOR2_X1 U557 ( .A(n738), .B(n737), .ZN(n767) );
  XNOR2_X1 U558 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n737) );
  XNOR2_X1 U559 ( .A(n780), .B(KEYINPUT105), .ZN(n782) );
  OR2_X1 U560 ( .A1(n832), .A2(n781), .ZN(n523) );
  INV_X1 U561 ( .A(KEYINPUT64), .ZN(n724) );
  NOR2_X1 U562 ( .A1(n717), .A2(n716), .ZN(n715) );
  XNOR2_X1 U563 ( .A(n775), .B(KEYINPUT32), .ZN(n776) );
  XNOR2_X1 U564 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X1 U565 ( .A1(n782), .A2(n523), .ZN(n783) );
  NOR2_X1 U566 ( .A1(n524), .A2(G2105), .ZN(n525) );
  INV_X1 U567 ( .A(KEYINPUT107), .ZN(n789) );
  XNOR2_X1 U568 ( .A(KEYINPUT72), .B(KEYINPUT13), .ZN(n591) );
  XNOR2_X1 U569 ( .A(n592), .B(n591), .ZN(n593) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n676) );
  XNOR2_X1 U571 ( .A(n539), .B(n538), .ZN(G160) );
  INV_X1 U572 ( .A(KEYINPUT65), .ZN(n539) );
  INV_X1 U573 ( .A(G2104), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT66), .ZN(n540) );
  NAND2_X1 U575 ( .A1(G101), .A2(n540), .ZN(n527) );
  INV_X1 U576 ( .A(KEYINPUT23), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n527), .B(n526), .ZN(n529) );
  AND2_X1 U578 ( .A1(n524), .A2(G2105), .ZN(n1004) );
  NAND2_X1 U579 ( .A1(n1004), .A2(G125), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X1 U581 ( .A(KEYINPUT67), .ZN(n530) );
  XNOR2_X1 U582 ( .A(n531), .B(n530), .ZN(n537) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT68), .B(n532), .Z(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT17), .B(n533), .ZN(n559) );
  NAND2_X1 U586 ( .A1(G137), .A2(n559), .ZN(n535) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n1005) );
  NAND2_X1 U588 ( .A1(n1005), .A2(G113), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U591 ( .A(n540), .ZN(n541) );
  INV_X1 U592 ( .A(n541), .ZN(n1008) );
  NAND2_X1 U593 ( .A1(G102), .A2(n1008), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G138), .A2(n559), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U596 ( .A1(G126), .A2(n1004), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G114), .A2(n1005), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U599 ( .A1(n547), .A2(n546), .ZN(G164) );
  XOR2_X1 U600 ( .A(G2454), .B(G2427), .Z(n549) );
  XNOR2_X1 U601 ( .A(G2451), .B(G2430), .ZN(n548) );
  XNOR2_X1 U602 ( .A(n549), .B(n548), .ZN(n556) );
  XOR2_X1 U603 ( .A(G2438), .B(G2435), .Z(n551) );
  XNOR2_X1 U604 ( .A(G1348), .B(G2446), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U606 ( .A(n552), .B(G2443), .Z(n554) );
  XNOR2_X1 U607 ( .A(G1341), .B(KEYINPUT109), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U610 ( .A1(n557), .A2(G14), .ZN(G401) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U612 ( .A1(G123), .A2(n1004), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n558), .B(KEYINPUT18), .ZN(n567) );
  NAND2_X1 U614 ( .A1(G99), .A2(n1008), .ZN(n562) );
  INV_X1 U615 ( .A(n559), .ZN(n560) );
  INV_X1 U616 ( .A(n560), .ZN(n1009) );
  NAND2_X1 U617 ( .A1(G135), .A2(n1009), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n1005), .A2(G111), .ZN(n563) );
  XOR2_X1 U620 ( .A(KEYINPUT80), .B(n563), .Z(n564) );
  NOR2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n1020) );
  XNOR2_X1 U623 ( .A(G2096), .B(n1020), .ZN(n568) );
  OR2_X1 U624 ( .A1(G2100), .A2(n568), .ZN(G156) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G82), .ZN(G220) );
  INV_X1 U627 ( .A(G96), .ZN(G221) );
  INV_X1 U628 ( .A(G120), .ZN(G236) );
  INV_X1 U629 ( .A(G69), .ZN(G235) );
  INV_X1 U630 ( .A(G108), .ZN(G238) );
  XOR2_X1 U631 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  INV_X1 U632 ( .A(G651), .ZN(n575) );
  NOR2_X1 U633 ( .A1(n649), .A2(n575), .ZN(n586) );
  NAND2_X1 U634 ( .A1(G76), .A2(n586), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G89), .A2(n676), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT4), .B(KEYINPUT78), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT79), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT5), .B(n574), .Z(n581) );
  NOR2_X1 U641 ( .A1(G543), .A2(n575), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT1), .B(n576), .Z(n672) );
  NAND2_X1 U643 ( .A1(G63), .A2(n672), .ZN(n578) );
  NOR2_X2 U644 ( .A1(G651), .A2(n649), .ZN(n675) );
  NAND2_X1 U645 ( .A1(G51), .A2(n675), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(KEYINPUT7), .B(n582), .ZN(G168) );
  XOR2_X1 U650 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n583) );
  XOR2_X1 U652 ( .A(n583), .B(KEYINPUT10), .Z(n1048) );
  NAND2_X1 U653 ( .A1(n1048), .A2(G567), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U655 ( .A1(n672), .A2(G56), .ZN(n585) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n585), .Z(n594) );
  NAND2_X1 U657 ( .A1(n586), .A2(G68), .ZN(n587) );
  XNOR2_X1 U658 ( .A(KEYINPUT71), .B(n587), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n676), .A2(G81), .ZN(n588) );
  XOR2_X1 U660 ( .A(n588), .B(KEYINPUT12), .Z(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n675), .A2(G43), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n1034) );
  INV_X1 U665 ( .A(G860), .ZN(n633) );
  OR2_X1 U666 ( .A1(n1034), .A2(n633), .ZN(G153) );
  NAND2_X1 U667 ( .A1(G77), .A2(n586), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G90), .A2(n676), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(KEYINPUT9), .B(n599), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G64), .A2(n672), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G52), .A2(n675), .ZN(n600) );
  AND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(G301) );
  INV_X1 U675 ( .A(G301), .ZN(G171) );
  INV_X1 U676 ( .A(G868), .ZN(n685) );
  NOR2_X1 U677 ( .A1(KEYINPUT73), .A2(G171), .ZN(n604) );
  NOR2_X1 U678 ( .A1(KEYINPUT77), .A2(n604), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n685), .A2(n605), .ZN(n621) );
  NAND2_X1 U680 ( .A1(G301), .A2(G868), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n606), .A2(KEYINPUT73), .ZN(n619) );
  NAND2_X1 U682 ( .A1(n675), .A2(G54), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n607), .Z(n609) );
  NAND2_X1 U684 ( .A1(n586), .A2(G79), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U686 ( .A(KEYINPUT76), .B(n610), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n672), .A2(G66), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT74), .B(n611), .Z(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n676), .A2(G92), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT15), .B(n616), .ZN(n1035) );
  NOR2_X1 U693 ( .A1(n1035), .A2(KEYINPUT77), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n685), .A2(n617), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n1035), .A2(KEYINPUT77), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(G284) );
  NAND2_X1 U699 ( .A1(G65), .A2(n672), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G78), .A2(n586), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n676), .A2(G91), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT70), .B(n626), .Z(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n675), .A2(G53), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(G299) );
  NOR2_X1 U707 ( .A1(G868), .A2(G299), .ZN(n632) );
  NOR2_X1 U708 ( .A1(G286), .A2(n685), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(G297) );
  NAND2_X1 U710 ( .A1(n633), .A2(G559), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n634), .A2(n1035), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U713 ( .A1(G868), .A2(n1034), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n1035), .A2(G868), .ZN(n636) );
  NOR2_X1 U715 ( .A1(G559), .A2(n636), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(G282) );
  NAND2_X1 U717 ( .A1(G75), .A2(n586), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G88), .A2(n676), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G62), .A2(n672), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G50), .A2(n675), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G49), .A2(n675), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U727 ( .A(KEYINPUT83), .B(n647), .Z(n648) );
  NOR2_X1 U728 ( .A1(n672), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G60), .A2(n672), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G72), .A2(n586), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G85), .A2(n676), .ZN(n654) );
  XNOR2_X1 U735 ( .A(KEYINPUT69), .B(n654), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n675), .A2(G47), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(G290) );
  NAND2_X1 U739 ( .A1(G61), .A2(n672), .ZN(n660) );
  NAND2_X1 U740 ( .A1(G86), .A2(n676), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n586), .A2(G73), .ZN(n661) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(n661), .Z(n662) );
  NOR2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n675), .A2(G48), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(G305) );
  NAND2_X1 U747 ( .A1(G559), .A2(n1035), .ZN(n666) );
  XOR2_X1 U748 ( .A(n1034), .B(n666), .Z(n975) );
  XOR2_X1 U749 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n668) );
  XNOR2_X1 U750 ( .A(G166), .B(KEYINPUT84), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n668), .B(n667), .ZN(n671) );
  XOR2_X1 U752 ( .A(G299), .B(G288), .Z(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(G290), .ZN(n670) );
  XNOR2_X1 U754 ( .A(n671), .B(n670), .ZN(n683) );
  NAND2_X1 U755 ( .A1(G67), .A2(n672), .ZN(n674) );
  NAND2_X1 U756 ( .A1(G80), .A2(n586), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n674), .A2(n673), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G55), .A2(n675), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G93), .A2(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U762 ( .A(KEYINPUT82), .B(n681), .Z(n978) );
  XNOR2_X1 U763 ( .A(G305), .B(n978), .ZN(n682) );
  XNOR2_X1 U764 ( .A(n683), .B(n682), .ZN(n1038) );
  XNOR2_X1 U765 ( .A(n975), .B(n1038), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n684), .A2(G868), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n685), .A2(n978), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n687), .A2(n686), .ZN(G295) );
  NAND2_X1 U769 ( .A1(G2084), .A2(G2078), .ZN(n688) );
  XOR2_X1 U770 ( .A(KEYINPUT20), .B(n688), .Z(n689) );
  NAND2_X1 U771 ( .A1(G2090), .A2(n689), .ZN(n690) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n690), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n691), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U774 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U775 ( .A1(G235), .A2(G236), .ZN(n692) );
  XNOR2_X1 U776 ( .A(n692), .B(KEYINPUT89), .ZN(n693) );
  NOR2_X1 U777 ( .A1(G238), .A2(n693), .ZN(n694) );
  NAND2_X1 U778 ( .A1(G57), .A2(n694), .ZN(n980) );
  NAND2_X1 U779 ( .A1(G567), .A2(n980), .ZN(n695) );
  XNOR2_X1 U780 ( .A(n695), .B(KEYINPUT90), .ZN(n703) );
  NOR2_X1 U781 ( .A1(G220), .A2(G219), .ZN(n696) );
  XOR2_X1 U782 ( .A(KEYINPUT22), .B(n696), .Z(n697) );
  NOR2_X1 U783 ( .A1(G218), .A2(n697), .ZN(n698) );
  XOR2_X1 U784 ( .A(KEYINPUT86), .B(n698), .Z(n699) );
  NOR2_X1 U785 ( .A1(G221), .A2(n699), .ZN(n700) );
  XNOR2_X1 U786 ( .A(KEYINPUT87), .B(n700), .ZN(n979) );
  NAND2_X1 U787 ( .A1(G2106), .A2(n979), .ZN(n701) );
  XNOR2_X1 U788 ( .A(KEYINPUT88), .B(n701), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U790 ( .A(n704), .B(KEYINPUT91), .Z(n981) );
  NAND2_X1 U791 ( .A1(G661), .A2(G483), .ZN(n705) );
  XNOR2_X1 U792 ( .A(KEYINPUT92), .B(n705), .ZN(n706) );
  NOR2_X1 U793 ( .A1(n981), .A2(n706), .ZN(n857) );
  NAND2_X1 U794 ( .A1(n857), .A2(G36), .ZN(G176) );
  XNOR2_X1 U795 ( .A(G166), .B(KEYINPUT93), .ZN(G303) );
  NOR2_X1 U796 ( .A1(G1976), .A2(G288), .ZN(n784) );
  NOR2_X1 U797 ( .A1(G1971), .A2(G303), .ZN(n707) );
  NOR2_X1 U798 ( .A1(n784), .A2(n707), .ZN(n959) );
  NOR2_X1 U799 ( .A1(G164), .A2(G1384), .ZN(n792) );
  AND2_X1 U800 ( .A1(G40), .A2(n792), .ZN(n708) );
  AND2_X1 U801 ( .A1(G160), .A2(n708), .ZN(n739) );
  INV_X1 U802 ( .A(n739), .ZN(n758) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n758), .ZN(n744) );
  NAND2_X1 U804 ( .A1(G8), .A2(n744), .ZN(n757) );
  NAND2_X1 U805 ( .A1(G8), .A2(n758), .ZN(n832) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n832), .ZN(n755) );
  INV_X1 U807 ( .A(G299), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G160), .A2(G40), .ZN(n791) );
  INV_X1 U809 ( .A(n792), .ZN(n710) );
  INV_X1 U810 ( .A(G2072), .ZN(n709) );
  OR2_X1 U811 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U812 ( .A1(n791), .A2(n711), .ZN(n712) );
  XNOR2_X1 U813 ( .A(n712), .B(KEYINPUT27), .ZN(n714) );
  AND2_X1 U814 ( .A1(G1956), .A2(n758), .ZN(n713) );
  NOR2_X1 U815 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U816 ( .A(n715), .B(KEYINPUT28), .Z(n731) );
  INV_X1 U817 ( .A(n731), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U819 ( .A1(n719), .A2(n718), .ZN(n736) );
  INV_X1 U820 ( .A(n1035), .ZN(n947) );
  AND2_X1 U821 ( .A1(n758), .A2(G1341), .ZN(n720) );
  OR2_X1 U822 ( .A1(n720), .A2(n1034), .ZN(n723) );
  INV_X1 U823 ( .A(G1996), .ZN(n992) );
  NOR2_X1 U824 ( .A1(n758), .A2(n992), .ZN(n721) );
  XNOR2_X1 U825 ( .A(n721), .B(KEYINPUT26), .ZN(n722) );
  NOR2_X1 U826 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U827 ( .A(n725), .B(n724), .ZN(n730) );
  OR2_X1 U828 ( .A1(n947), .A2(n730), .ZN(n729) );
  NOR2_X1 U829 ( .A1(G2067), .A2(n758), .ZN(n727) );
  NOR2_X1 U830 ( .A1(n739), .A2(G1348), .ZN(n726) );
  NOR2_X1 U831 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U832 ( .A1(n729), .A2(n728), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n730), .A2(n947), .ZN(n732) );
  AND2_X1 U834 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U836 ( .A1(n736), .A2(n735), .ZN(n738) );
  INV_X1 U837 ( .A(G1961), .ZN(n985) );
  NAND2_X1 U838 ( .A1(n758), .A2(n985), .ZN(n741) );
  XNOR2_X1 U839 ( .A(G2078), .B(KEYINPUT25), .ZN(n899) );
  NAND2_X1 U840 ( .A1(n739), .A2(n899), .ZN(n740) );
  NAND2_X1 U841 ( .A1(n741), .A2(n740), .ZN(n743) );
  AND2_X1 U842 ( .A1(n743), .A2(G171), .ZN(n742) );
  XOR2_X1 U843 ( .A(KEYINPUT98), .B(n742), .Z(n765) );
  NAND2_X1 U844 ( .A1(n767), .A2(n765), .ZN(n752) );
  NOR2_X1 U845 ( .A1(G171), .A2(n743), .ZN(n749) );
  NOR2_X1 U846 ( .A1(n755), .A2(n744), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U848 ( .A(n746), .B(KEYINPUT30), .ZN(n747) );
  NOR2_X1 U849 ( .A1(G168), .A2(n747), .ZN(n748) );
  NOR2_X1 U850 ( .A1(n749), .A2(n748), .ZN(n751) );
  XOR2_X1 U851 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n750) );
  XNOR2_X1 U852 ( .A(n751), .B(n750), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n752), .A2(n770), .ZN(n753) );
  XNOR2_X1 U854 ( .A(n753), .B(KEYINPUT101), .ZN(n754) );
  NOR2_X1 U855 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U856 ( .A1(n757), .A2(n756), .ZN(n779) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n832), .ZN(n760) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U859 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U860 ( .A1(n761), .A2(G303), .ZN(n762) );
  XNOR2_X1 U861 ( .A(n762), .B(KEYINPUT102), .ZN(n769) );
  INV_X1 U862 ( .A(n769), .ZN(n763) );
  OR2_X1 U863 ( .A1(n763), .A2(G286), .ZN(n764) );
  AND2_X1 U864 ( .A1(n764), .A2(G8), .ZN(n768) );
  AND2_X1 U865 ( .A1(n765), .A2(n768), .ZN(n766) );
  NAND2_X1 U866 ( .A1(n767), .A2(n766), .ZN(n774) );
  INV_X1 U867 ( .A(n768), .ZN(n772) );
  AND2_X1 U868 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  AND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n777) );
  XOR2_X1 U871 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n775) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n828) );
  NAND2_X1 U873 ( .A1(n959), .A2(n828), .ZN(n780) );
  NAND2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NOR2_X1 U875 ( .A1(KEYINPUT33), .A2(n783), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n784), .A2(KEYINPUT33), .ZN(n785) );
  XNOR2_X1 U877 ( .A(KEYINPUT106), .B(n785), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n786), .A2(n832), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n790), .B(n789), .ZN(n823) );
  XOR2_X1 U881 ( .A(G1981), .B(G305), .Z(n952) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n848) );
  XNOR2_X1 U883 ( .A(G1986), .B(G290), .ZN(n964) );
  NAND2_X1 U884 ( .A1(n848), .A2(n964), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT94), .B(n793), .ZN(n825) );
  AND2_X1 U886 ( .A1(n952), .A2(n825), .ZN(n821) );
  NAND2_X1 U887 ( .A1(n1005), .A2(G107), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G95), .A2(n1008), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G119), .A2(n1004), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G131), .A2(n1009), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n1027) );
  XOR2_X1 U894 ( .A(G1991), .B(KEYINPUT97), .Z(n900) );
  AND2_X1 U895 ( .A1(n1027), .A2(n900), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G129), .A2(n1004), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G141), .A2(n1009), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G105), .A2(n1008), .ZN(n802) );
  XNOR2_X1 U900 ( .A(n802), .B(KEYINPUT38), .ZN(n804) );
  NAND2_X1 U901 ( .A1(G117), .A2(n1005), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n1021) );
  NOR2_X1 U904 ( .A1(n992), .A2(n1021), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n840) );
  NAND2_X1 U906 ( .A1(G128), .A2(n1004), .ZN(n810) );
  NAND2_X1 U907 ( .A1(G116), .A2(n1005), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U909 ( .A(KEYINPUT35), .B(n811), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G140), .A2(n1009), .ZN(n812) );
  XNOR2_X1 U911 ( .A(n812), .B(KEYINPUT96), .ZN(n814) );
  NAND2_X1 U912 ( .A1(G104), .A2(n1008), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U914 ( .A(KEYINPUT34), .B(n815), .Z(n816) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U916 ( .A(KEYINPUT36), .B(n818), .Z(n1030) );
  XNOR2_X1 U917 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  XOR2_X1 U918 ( .A(n819), .B(KEYINPUT95), .Z(n839) );
  OR2_X1 U919 ( .A1(n1030), .A2(n839), .ZN(n889) );
  NAND2_X1 U920 ( .A1(n840), .A2(n889), .ZN(n820) );
  NAND2_X1 U921 ( .A1(n820), .A2(n848), .ZN(n824) );
  AND2_X1 U922 ( .A1(n821), .A2(n824), .ZN(n822) );
  NAND2_X1 U923 ( .A1(n823), .A2(n822), .ZN(n853) );
  INV_X1 U924 ( .A(n824), .ZN(n838) );
  INV_X1 U925 ( .A(n825), .ZN(n836) );
  NOR2_X1 U926 ( .A1(G2090), .A2(G303), .ZN(n826) );
  NAND2_X1 U927 ( .A1(G8), .A2(n826), .ZN(n827) );
  NAND2_X1 U928 ( .A1(n828), .A2(n827), .ZN(n829) );
  AND2_X1 U929 ( .A1(n829), .A2(n832), .ZN(n834) );
  NOR2_X1 U930 ( .A1(G1981), .A2(G305), .ZN(n830) );
  XOR2_X1 U931 ( .A(n830), .B(KEYINPUT24), .Z(n831) );
  NOR2_X1 U932 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n835) );
  OR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  OR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n851) );
  NAND2_X1 U936 ( .A1(n1030), .A2(n839), .ZN(n888) );
  AND2_X1 U937 ( .A1(n992), .A2(n1021), .ZN(n876) );
  INV_X1 U938 ( .A(n840), .ZN(n881) );
  NOR2_X1 U939 ( .A1(G1986), .A2(G290), .ZN(n841) );
  NOR2_X1 U940 ( .A1(n900), .A2(n1027), .ZN(n884) );
  NOR2_X1 U941 ( .A1(n841), .A2(n884), .ZN(n842) );
  NOR2_X1 U942 ( .A1(n881), .A2(n842), .ZN(n843) );
  NOR2_X1 U943 ( .A1(n876), .A2(n843), .ZN(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT39), .B(n844), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT108), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n846), .A2(n889), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n888), .A2(n847), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n850) );
  AND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U950 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U952 ( .A1(G2106), .A2(n1048), .ZN(G217) );
  AND2_X1 U953 ( .A1(G15), .A2(G2), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G661), .A2(n855), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(G188) );
  NAND2_X1 U958 ( .A1(n1004), .A2(G124), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G112), .A2(n1005), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G100), .A2(n1008), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G136), .A2(n1009), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(G162) );
  INV_X1 U966 ( .A(KEYINPUT55), .ZN(n894) );
  NAND2_X1 U967 ( .A1(G103), .A2(n1008), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G139), .A2(n1009), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G127), .A2(n1004), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G115), .A2(n1005), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n1026) );
  XOR2_X1 U975 ( .A(G2072), .B(n1026), .Z(n873) );
  XOR2_X1 U976 ( .A(G164), .B(G2078), .Z(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U978 ( .A(KEYINPUT50), .B(n874), .ZN(n879) );
  XOR2_X1 U979 ( .A(G2090), .B(G162), .Z(n875) );
  NOR2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(KEYINPUT51), .B(n877), .Z(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n887) );
  XNOR2_X1 U984 ( .A(G160), .B(G2084), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n882), .A2(n1020), .ZN(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(KEYINPUT118), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(KEYINPUT52), .B(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n895), .A2(G29), .ZN(n945) );
  XNOR2_X1 U994 ( .A(G2090), .B(G35), .ZN(n910) );
  XOR2_X1 U995 ( .A(G32), .B(G1996), .Z(n896) );
  NAND2_X1 U996 ( .A1(n896), .A2(G28), .ZN(n906) );
  XNOR2_X1 U997 ( .A(G2067), .B(G26), .ZN(n898) );
  XNOR2_X1 U998 ( .A(G33), .B(G2072), .ZN(n897) );
  NOR2_X1 U999 ( .A1(n898), .A2(n897), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n899), .B(G27), .Z(n902) );
  XNOR2_X1 U1001 ( .A(n900), .B(G25), .ZN(n901) );
  NOR2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT119), .B(n907), .Z(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT53), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G2084), .B(KEYINPUT54), .Z(n911) );
  XNOR2_X1 U1009 ( .A(G34), .B(n911), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(KEYINPUT55), .B(n914), .Z(n916) );
  INV_X1 U1012 ( .A(G29), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(G11), .A2(n917), .ZN(n943) );
  XOR2_X1 U1015 ( .A(G20), .B(G1956), .Z(n921) );
  XNOR2_X1 U1016 ( .A(G1341), .B(G19), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1021 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT60), .B(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(G1961), .B(G5), .Z(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G21), .B(G1966), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT124), .B(n930), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G1976), .B(G23), .Z(n932) );
  XOR2_X1 U1030 ( .A(G1971), .B(G22), .Z(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G24), .B(G1986), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(n938), .B(KEYINPUT61), .Z(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT125), .B(n939), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n940), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(KEYINPUT126), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n973) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .Z(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n946), .ZN(n971) );
  XOR2_X1 U1044 ( .A(G1348), .B(n947), .Z(n951) );
  XOR2_X1 U1045 ( .A(G171), .B(G1961), .Z(n949) );
  XNOR2_X1 U1046 ( .A(n1034), .B(G1341), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n969) );
  XNOR2_X1 U1049 ( .A(G168), .B(G1966), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT121), .ZN(n955) );
  XOR2_X1 U1052 ( .A(KEYINPUT57), .B(n955), .Z(n967) );
  XOR2_X1 U1053 ( .A(G299), .B(G1956), .Z(n957) );
  NAND2_X1 U1054 ( .A1(G1971), .A2(G303), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT122), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1060 ( .A(KEYINPUT123), .B(n965), .Z(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n974), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1066 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  XNOR2_X1 U1067 ( .A(n975), .B(KEYINPUT81), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(G860), .A2(n976), .ZN(n977) );
  XOR2_X1 U1069 ( .A(n978), .B(n977), .Z(G145) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(G325) );
  INV_X1 U1071 ( .A(G325), .ZN(G261) );
  INV_X1 U1072 ( .A(n981), .ZN(G319) );
  XOR2_X1 U1073 ( .A(KEYINPUT111), .B(G2474), .Z(n983) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G1976), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1076 ( .A(n984), .B(KEYINPUT41), .Z(n987) );
  XOR2_X1 U1077 ( .A(n985), .B(G1956), .Z(n986) );
  XNOR2_X1 U1078 ( .A(n987), .B(n986), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT112), .B(G1986), .Z(n989) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G1971), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n989), .B(n988), .ZN(n990) );
  XOR2_X1 U1082 ( .A(n991), .B(n990), .Z(n994) );
  XOR2_X1 U1083 ( .A(n992), .B(G1991), .Z(n993) );
  XNOR2_X1 U1084 ( .A(n994), .B(n993), .ZN(G229) );
  XOR2_X1 U1085 ( .A(G2100), .B(G2096), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G2090), .B(KEYINPUT43), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n996), .B(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(n997), .B(KEYINPUT110), .Z(n999) );
  XNOR2_X1 U1089 ( .A(G2072), .B(G2678), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n999), .B(n998), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT42), .B(G2067), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(G2084), .B(G2078), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1003), .B(n1002), .ZN(G227) );
  NAND2_X1 U1095 ( .A1(G130), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(G118), .A2(n1005), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(G106), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(G142), .A2(n1009), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT45), .B(n1012), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT114), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT113), .B(KEYINPUT115), .Z(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1019), .B(n1018), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(n1020), .B(G162), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(G164), .B(n1021), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(n1023), .B(n1022), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(n1025), .B(n1024), .Z(n1029) );
  XOR2_X1 U1112 ( .A(n1027), .B(n1026), .Z(n1028) );
  XNOR2_X1 U1113 ( .A(n1029), .B(n1028), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(n1030), .B(G160), .Z(n1031) );
  XNOR2_X1 U1115 ( .A(n1032), .B(n1031), .ZN(n1033) );
  NOR2_X1 U1116 ( .A1(G37), .A2(n1033), .ZN(G395) );
  XNOR2_X1 U1117 ( .A(n1034), .B(KEYINPUT116), .ZN(n1037) );
  XOR2_X1 U1118 ( .A(G301), .B(n1035), .Z(n1036) );
  XNOR2_X1 U1119 ( .A(n1037), .B(n1036), .ZN(n1040) );
  XNOR2_X1 U1120 ( .A(G286), .B(n1038), .ZN(n1039) );
  XNOR2_X1 U1121 ( .A(n1040), .B(n1039), .ZN(n1041) );
  NOR2_X1 U1122 ( .A1(G37), .A2(n1041), .ZN(G397) );
  NOR2_X1 U1123 ( .A1(G229), .A2(G227), .ZN(n1042) );
  XNOR2_X1 U1124 ( .A(n1042), .B(KEYINPUT49), .ZN(n1043) );
  NOR2_X1 U1125 ( .A1(G401), .A2(n1043), .ZN(n1044) );
  NAND2_X1 U1126 ( .A1(G319), .A2(n1044), .ZN(n1045) );
  XNOR2_X1 U1127 ( .A(KEYINPUT117), .B(n1045), .ZN(n1047) );
  NOR2_X1 U1128 ( .A1(G395), .A2(G397), .ZN(n1046) );
  NAND2_X1 U1129 ( .A1(n1047), .A2(n1046), .ZN(G225) );
  INV_X1 U1130 ( .A(G225), .ZN(G308) );
  INV_X1 U1131 ( .A(G57), .ZN(G237) );
  INV_X1 U1132 ( .A(n1048), .ZN(G223) );
endmodule

