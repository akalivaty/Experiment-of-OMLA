//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n189), .A2(new_n192), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n188), .A2(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT68), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT68), .A2(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(G116), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT5), .A3(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT68), .A2(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT68), .A2(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT5), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G116), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(G113), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n212));
  INV_X1    g026(.A(new_n204), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(new_n208), .B2(G116), .ZN(new_n214));
  INV_X1    g028(.A(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n212), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n212), .A2(new_n202), .A3(new_n204), .A4(new_n219), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n199), .B(new_n211), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n202), .A2(new_n204), .ZN(new_n223));
  INV_X1    g037(.A(new_n219), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n212), .A3(new_n219), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n225), .A2(new_n226), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n189), .A2(new_n192), .A3(new_n194), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n195), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n222), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n187), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n222), .B(new_n235), .C1(new_n227), .C2(new_n233), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n187), .A3(new_n236), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n234), .A2(KEYINPUT81), .A3(new_n187), .A4(new_n236), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT0), .A3(G128), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(G143), .B(G146), .Z(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n256), .B(G128), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G128), .B1(new_n259), .B2(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n254), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(KEYINPUT82), .A3(G125), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n255), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT83), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n242), .A2(new_n247), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n238), .B(new_n239), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n274), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n255), .A2(new_n264), .A3(new_n265), .A4(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n211), .B1(new_n220), .B2(new_n221), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n195), .A2(new_n198), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n222), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n235), .B(KEYINPUT8), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n275), .A2(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n272), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n286), .B(KEYINPUT84), .Z(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n286), .A3(new_n284), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT85), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n287), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT85), .B(new_n291), .C1(new_n271), .C2(new_n284), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G214), .B1(G237), .B2(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G140), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT77), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n267), .A2(G227), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n233), .B2(new_n252), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n253), .A2(new_n230), .A3(KEYINPUT78), .A4(new_n232), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G137), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT64), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G137), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT11), .A2(G134), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT65), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(G134), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n310), .A2(new_n312), .A3(new_n313), .A4(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G134), .ZN(new_n321));
  AOI21_X1  g135(.A(G131), .B1(new_n321), .B2(G137), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n315), .A2(new_n318), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT66), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n320), .A2(new_n318), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n315), .A4(new_n322), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(G137), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n315), .A2(new_n318), .A3(new_n320), .A4(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n324), .A2(new_n327), .B1(G131), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n199), .A2(new_n262), .A3(new_n260), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT10), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n199), .A2(new_n333), .A3(new_n262), .A4(new_n260), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n308), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n306), .A2(new_n307), .B1(new_n334), .B2(new_n332), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n330), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n304), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n263), .A2(new_n279), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n331), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(new_n330), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n324), .A2(new_n327), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n329), .A2(G131), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n343), .A3(KEYINPUT12), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n336), .A3(new_n303), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n345), .A2(new_n349), .B1(new_n338), .B2(new_n330), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n336), .A2(new_n303), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n356), .A2(new_n303), .B1(new_n357), .B2(new_n339), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n359), .B2(KEYINPUT79), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n361), .B(new_n353), .C1(new_n358), .C2(new_n354), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n297), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G478), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT15), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n296), .A2(new_n367), .A3(G953), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G128), .B(G143), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(new_n321), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  INV_X1    g186(.A(G122), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G116), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n203), .A2(KEYINPUT92), .A3(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n203), .B2(G122), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n371), .B1(G107), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n374), .B2(new_n375), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n380), .A2(new_n381), .B1(G116), .B2(new_n373), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n374), .A2(new_n375), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT93), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT94), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n379), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n378), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(G134), .C1(new_n258), .C2(G128), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n371), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n377), .B(new_n191), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n369), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n385), .A2(KEYINPUT94), .B1(new_n379), .B2(new_n383), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n191), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n398), .B(new_n368), .C1(new_n400), .C2(new_n378), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n366), .B1(new_n402), .B2(new_n354), .ZN(new_n403));
  AOI211_X1 g217(.A(G902), .B(new_n365), .C1(new_n397), .C2(new_n401), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n354), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT21), .B(G898), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR2_X1    g221(.A1(KEYINPUT95), .A2(G952), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT95), .A2(G952), .ZN(new_n409));
  AOI21_X1  g223(.A(G953), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G234), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n403), .A2(new_n404), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  NOR2_X1   g231(.A1(G237), .A2(G953), .ZN(new_n418));
  AOI21_X1  g232(.A(G143), .B1(new_n418), .B2(G214), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(G143), .A3(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  INV_X1    g238(.A(G131), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n425), .A3(new_n421), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n254), .A2(KEYINPUT72), .A3(G140), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G125), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n254), .A2(G140), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT72), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(KEYINPUT16), .ZN(new_n434));
  INV_X1    g248(.A(G146), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT16), .B1(new_n430), .B2(G125), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G146), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n427), .A2(new_n438), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G125), .B(G140), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n428), .B1(new_n443), .B2(KEYINPUT72), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G146), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n435), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT18), .A2(G131), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n420), .A2(new_n421), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n422), .A2(KEYINPUT18), .A3(G131), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT87), .B(G104), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT89), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n454), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n442), .B2(new_n451), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n354), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n417), .B1(new_n460), .B2(KEYINPUT91), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(new_n354), .C1(new_n457), .C2(new_n459), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n436), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(new_n435), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n439), .A2(KEYINPUT73), .A3(G146), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n423), .A2(new_n426), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n443), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n429), .A2(new_n433), .B1(new_n443), .B2(KEYINPUT86), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n435), .B(new_n472), .C1(new_n473), .C2(new_n471), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n458), .B1(new_n475), .B2(new_n451), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI211_X1 g292(.A(KEYINPUT88), .B(new_n458), .C1(new_n475), .C2(new_n451), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n456), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n481), .A2(new_n482), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n485), .A3(new_n482), .A4(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n416), .B(new_n464), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n295), .A2(new_n363), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  INV_X1    g304(.A(new_n316), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n310), .A2(new_n312), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(new_n321), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n260), .B(new_n262), .C1(new_n493), .C2(new_n425), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n327), .B2(new_n324), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n348), .B2(new_n253), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n496), .B2(new_n227), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n346), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n330), .B2(new_n252), .ZN(new_n501));
  INV_X1    g315(.A(new_n227), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n418), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G101), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT29), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n501), .A2(KEYINPUT28), .A3(new_n502), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n507), .B1(new_n515), .B2(new_n497), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT70), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n517), .A3(new_n354), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n348), .A2(new_n519), .A3(new_n253), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT67), .B1(new_n330), .B2(new_n252), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n495), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI22_X1  g336(.A1(new_n515), .A2(new_n497), .B1(new_n522), .B2(new_n227), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n511), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n503), .A2(new_n511), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n522), .A2(KEYINPUT30), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n500), .B(KEYINPUT30), .C1(new_n330), .C2(new_n252), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n502), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n525), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G472), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n519), .B1(new_n348), .B2(new_n253), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n330), .A2(KEYINPUT67), .A3(new_n252), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n500), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n496), .A2(new_n227), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n511), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT31), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n511), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n523), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n503), .A2(new_n540), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n542), .B(new_n543), .C1(new_n526), .C2(new_n528), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n531), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n367), .B1(G234), .B2(new_n354), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  INV_X1    g371(.A(G128), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT23), .A3(G119), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT71), .B(new_n558), .C1(new_n206), .C2(new_n207), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n206), .A2(new_n207), .A3(new_n558), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n200), .A2(new_n201), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT71), .B1(new_n564), .B2(new_n558), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n557), .B(new_n559), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n558), .A2(G119), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n564), .B2(new_n558), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT24), .B(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n467), .A3(new_n468), .A4(new_n446), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n440), .A2(new_n438), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n559), .B1(new_n563), .B2(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G110), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n568), .A2(new_n569), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n572), .A2(KEYINPUT74), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT74), .B1(new_n572), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n556), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n577), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n555), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT25), .B1(new_n583), .B2(new_n354), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n585), .B(G902), .C1(new_n580), .C2(new_n582), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n551), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n582), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n572), .A2(new_n577), .A3(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n592), .B2(new_n556), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n551), .A2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n587), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n489), .A2(new_n550), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n545), .A2(new_n354), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n545), .A2(new_n547), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n363), .A2(new_n596), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n464), .B1(new_n484), .B2(new_n487), .ZN(new_n605));
  INV_X1    g419(.A(new_n294), .ZN(new_n606));
  INV_X1    g420(.A(new_n286), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n285), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n608), .B2(new_n289), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT33), .B1(new_n368), .B2(KEYINPUT96), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n402), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n397), .A2(new_n401), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n364), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n402), .A2(new_n354), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(G478), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n364), .A2(new_n354), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n605), .A2(new_n609), .A3(new_n618), .A4(new_n414), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n603), .A2(new_n604), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n403), .ZN(new_n623));
  INV_X1    g437(.A(new_n404), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n414), .B(KEYINPUT97), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n464), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n271), .A2(new_n286), .A3(new_n284), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n286), .B1(new_n271), .B2(new_n284), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n294), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n480), .A2(new_n483), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n482), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n480), .A2(KEYINPUT20), .A3(new_n483), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n603), .A2(new_n604), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n555), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n578), .B2(new_n579), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n640), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n590), .A2(new_n591), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT99), .B1(new_n646), .B2(new_n594), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n648), .B(new_n595), .C1(new_n642), .C2(new_n645), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n587), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n601), .A2(new_n602), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n601), .A2(new_n654), .A3(new_n651), .A4(new_n602), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n489), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n551), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n585), .B1(new_n593), .B2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n583), .A2(KEYINPUT25), .A3(new_n354), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n578), .A2(new_n641), .A3(new_n579), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n644), .B1(new_n590), .B2(new_n591), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n594), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n648), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n646), .A2(KEYINPUT99), .A3(new_n594), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n363), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n403), .A2(new_n404), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n405), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n673), .A2(new_n413), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n461), .B2(new_n463), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n632), .A2(new_n675), .A3(new_n633), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n630), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n550), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NAND2_X1  g493(.A1(new_n290), .A2(new_n293), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n605), .A2(new_n625), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n606), .A3(new_n651), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n511), .B1(new_n536), .B2(new_n503), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n525), .ZN(new_n687));
  INV_X1    g501(.A(new_n507), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n354), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n548), .B2(new_n549), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n682), .A2(new_n684), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n682), .A2(new_n684), .A3(new_n694), .A4(new_n691), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n674), .B(KEYINPUT39), .Z(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n363), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT40), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n693), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n693), .A2(new_n702), .A3(new_n695), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n258), .ZN(G45));
  INV_X1    g519(.A(new_n674), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n605), .A2(new_n609), .A3(new_n618), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n670), .A2(new_n707), .A3(new_n550), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  AOI21_X1  g523(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n297), .A3(new_n355), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n596), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n619), .A2(new_n550), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n550), .A2(new_n713), .A3(new_n635), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR2_X1   g532(.A1(new_n669), .A2(new_n488), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n630), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n550), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT104), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n719), .A2(new_n550), .A3(new_n723), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND2_X1  g540(.A1(new_n475), .A2(new_n451), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n454), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT88), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n476), .A2(new_n477), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n457), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n482), .B1(new_n731), .B2(new_n485), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n631), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n733), .A2(new_n486), .B1(new_n463), .B2(new_n461), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n630), .A3(new_n671), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n516), .A2(new_n540), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n539), .A2(new_n544), .A3(new_n736), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n600), .A2(G472), .B1(new_n547), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n626), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n712), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n597), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  AND3_X1   g556(.A1(new_n605), .A2(new_n618), .A3(new_n706), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n720), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n737), .A2(new_n547), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n601), .A2(new_n651), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n651), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n254), .ZN(G27));
  XOR2_X1   g565(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n550), .A2(new_n597), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n606), .B1(new_n290), .B2(new_n293), .ZN(new_n755));
  INV_X1    g569(.A(new_n297), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n357), .A2(new_n339), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n303), .B1(new_n350), .B2(new_n336), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n759), .B2(G902), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n760), .B2(new_n355), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n743), .A2(new_n755), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n753), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n680), .A2(new_n294), .A3(new_n761), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n605), .A2(new_n618), .A3(new_n706), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n550), .A3(new_n597), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n676), .A2(new_n671), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n755), .A2(new_n773), .A3(new_n761), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n754), .B2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n755), .A2(new_n773), .A3(new_n761), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n550), .A4(new_n597), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  NAND2_X1  g593(.A1(new_n734), .A2(new_n618), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT43), .Z(new_n781));
  NOR2_X1   g595(.A1(new_n603), .A2(new_n669), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT44), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n759), .A2(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(G469), .B1(new_n759), .B2(KEYINPUT45), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(G469), .A2(G902), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n787), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n355), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n297), .A3(new_n696), .ZN(new_n793));
  INV_X1    g607(.A(new_n755), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n783), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT108), .B(G137), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  NAND2_X1  g613(.A1(new_n792), .A2(new_n297), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n297), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n550), .A2(new_n794), .A3(new_n597), .A4(new_n765), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  INV_X1    g621(.A(new_n413), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n781), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n597), .A2(new_n738), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n355), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n710), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n816), .A2(new_n756), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n755), .B1(new_n804), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n606), .B1(new_n820), .B2(KEYINPUT50), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n682), .A2(new_n712), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n812), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n809), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n794), .A2(new_n712), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT105), .B1(new_n738), .B2(new_n651), .ZN(new_n829));
  AND4_X1   g643(.A1(KEYINPUT105), .A2(new_n601), .A3(new_n651), .A4(new_n745), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n691), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n597), .A3(new_n832), .A4(new_n808), .ZN(new_n833));
  OR3_X1    g647(.A1(new_n833), .A2(new_n605), .A3(new_n618), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n823), .B1(new_n811), .B2(new_n822), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n837), .ZN(new_n841));
  INV_X1    g655(.A(new_n754), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n842), .A3(new_n828), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n605), .A2(new_n618), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n814), .A2(new_n609), .A3(new_n297), .ZN(new_n847));
  OAI221_X1 g661(.A(new_n410), .B1(new_n846), .B2(new_n833), .C1(new_n812), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n840), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n775), .A2(new_n777), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT109), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT109), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n403), .B2(new_n404), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n734), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n846), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n295), .A2(new_n739), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n603), .A2(new_n857), .A3(new_n604), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n656), .A2(new_n598), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n766), .B1(new_n830), .B2(new_n829), .ZN(new_n861));
  INV_X1    g675(.A(new_n676), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT110), .A3(new_n852), .A4(new_n854), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(new_n755), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n855), .B2(new_n676), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n550), .A3(new_n670), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n851), .A2(new_n860), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n550), .B(new_n670), .C1(new_n707), .C2(new_n677), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n605), .A2(new_n761), .A3(new_n609), .A4(new_n625), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n651), .B2(new_n674), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n587), .A2(new_n650), .A3(KEYINPUT111), .A4(new_n706), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n871), .A2(new_n691), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT112), .B1(new_n876), .B2(new_n750), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n847), .A2(new_n765), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n830), .B2(new_n829), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n870), .A4(new_n875), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n714), .A2(new_n717), .A3(new_n741), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n770), .A2(new_n725), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n869), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT52), .B1(new_n877), .B2(new_n881), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT53), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(new_n876), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n879), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n877), .A2(new_n881), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n888), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n884), .A4(new_n869), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n887), .A2(new_n894), .A3(KEYINPUT54), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n885), .B2(new_n886), .ZN(new_n896));
  INV_X1    g710(.A(new_n868), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n656), .A2(new_n598), .A3(new_n859), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n778), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT113), .A4(new_n778), .ZN(new_n902));
  INV_X1    g716(.A(new_n770), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n725), .A2(new_n883), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n893), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n892), .A2(new_n901), .A3(new_n902), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n896), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n895), .A2(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n850), .A2(new_n909), .B1(G952), .B2(G953), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n756), .B(new_n606), .C1(new_n815), .C2(KEYINPUT49), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT49), .B2(new_n815), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n596), .A3(new_n780), .ZN(new_n913));
  INV_X1    g727(.A(new_n682), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n832), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(G75));
  OR2_X1    g730(.A1(new_n267), .A2(G952), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT118), .Z(new_n918));
  AOI211_X1 g732(.A(new_n354), .B(new_n291), .C1(new_n896), .C2(new_n906), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n242), .A2(new_n247), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n270), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT55), .Z(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n354), .B1(new_n896), .B2(new_n906), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  INV_X1    g741(.A(new_n922), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(G210), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n930), .B(new_n354), .C1(new_n896), .C2(new_n906), .ZN(new_n931));
  OAI211_X1 g745(.A(KEYINPUT117), .B(new_n922), .C1(new_n931), .C2(KEYINPUT56), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n929), .B2(new_n932), .ZN(G51));
  INV_X1    g747(.A(new_n918), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n787), .B(KEYINPUT57), .Z(new_n935));
  INV_X1    g749(.A(new_n908), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n907), .B1(new_n896), .B2(new_n906), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n352), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n786), .B(KEYINPUT119), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n926), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n934), .B1(new_n939), .B2(new_n941), .ZN(G54));
  NAND3_X1  g756(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(new_n480), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n480), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n934), .B1(new_n944), .B2(new_n945), .ZN(G60));
  NAND2_X1  g760(.A1(new_n611), .A2(new_n613), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT120), .Z(new_n948));
  XOR2_X1   g762(.A(new_n617), .B(KEYINPUT59), .Z(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n949), .C1(new_n936), .C2(new_n937), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n918), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n909), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(new_n896), .A2(new_n906), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n367), .A2(new_n354), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n934), .B1(new_n958), .B2(new_n593), .ZN(new_n959));
  INV_X1    g773(.A(new_n957), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n896), .B2(new_n906), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n646), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n959), .B(new_n962), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT122), .B(new_n918), .C1(new_n961), .C2(new_n583), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n918), .B1(new_n961), .B2(new_n583), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n954), .A2(new_n646), .A3(new_n957), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n406), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n267), .B1(new_n970), .B2(G224), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n904), .A2(new_n860), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(new_n267), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n920), .B1(G898), .B2(new_n267), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(G69));
  AOI21_X1  g790(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n842), .A2(new_n698), .A3(new_n755), .A4(new_n857), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT125), .Z(new_n979));
  NAND3_X1  g793(.A1(new_n797), .A2(new_n979), .A3(new_n806), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n879), .A2(new_n870), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n701), .A2(new_n703), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n701), .A2(KEYINPUT62), .A3(new_n703), .A4(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n527), .B1(new_n522), .B2(KEYINPUT30), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT123), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT124), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n851), .B1(new_n795), .B2(new_n796), .ZN(new_n994));
  NOR4_X1   g808(.A1(new_n793), .A2(new_n754), .A3(new_n630), .A4(new_n683), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n804), .B2(new_n805), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n994), .A2(new_n996), .A3(new_n770), .A4(new_n981), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(G953), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n672), .B2(new_n267), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n977), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n977), .ZN(new_n1002));
  OAI221_X1 g816(.A(new_n1002), .B1(new_n998), .B2(new_n999), .C1(new_n987), .C2(new_n992), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  AND3_X1   g820(.A1(new_n685), .A2(new_n529), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n887), .A2(new_n894), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n997), .A2(new_n973), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1006), .B(KEYINPUT126), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n918), .B(new_n1008), .C1(new_n1012), .C2(new_n529), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n986), .B2(new_n972), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n685), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(G57));
endmodule


