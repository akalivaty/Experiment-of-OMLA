//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1189, new_n1190, new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n477), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n477), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n467), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(KEYINPUT70), .A3(G138), .A4(new_n477), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n485), .A2(new_n486), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n509), .A3(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n502), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AND3_X1   g091(.A1(new_n507), .A2(new_n509), .A3(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G51), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n499), .A2(G89), .A3(new_n507), .A4(new_n509), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n504), .A2(new_n506), .A3(G63), .A4(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n510), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n519), .A2(new_n521), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n512), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT71), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G52), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n510), .A2(new_n534), .B1(new_n536), .B2(new_n512), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n499), .B2(G64), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n501), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n504), .A2(new_n506), .A3(G64), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n537), .B1(new_n542), .B2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n501), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n510), .A2(new_n549), .B1(new_n512), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  AOI22_X1  g134(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n501), .B1(new_n561), .B2(new_n510), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n507), .A2(new_n509), .A3(G53), .A4(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  AND4_X1   g142(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G90), .B1(new_n517), .B2(new_n535), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n543), .A2(new_n541), .A3(new_n538), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n541), .B1(new_n543), .B2(new_n538), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n568), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n517), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  AOI22_X1  g153(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n501), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n510), .A2(new_n581), .B1(new_n512), .B2(new_n582), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n580), .A2(new_n583), .A3(KEYINPUT75), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT75), .B1(new_n580), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G305));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n510), .A2(new_n587), .B1(new_n512), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n590), .A2(new_n591), .B1(new_n501), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n499), .A2(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n510), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G299), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n552), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n613), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n617), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n620), .B1(new_n623), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n493), .A2(new_n469), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n478), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n468), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n477), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n657), .B2(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n660), .B1(new_n659), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n671));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n668), .A2(new_n669), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(new_n681), .B(new_n680), .S(new_n673), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT85), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n683), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(new_n469), .A2(G103), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT25), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G139), .ZN(new_n695));
  INV_X1    g270(.A(new_n468), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(new_n477), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G33), .B(new_n701), .S(G29), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G2072), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G171), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G5), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT95), .B(G1961), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT29), .Z(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n709), .B1(KEYINPUT24), .B2(G34), .ZN(new_n716));
  OAI22_X1  g291(.A1(G160), .A2(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2084), .ZN(new_n718));
  NOR2_X1   g293(.A1(G29), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n478), .A2(G129), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n468), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n469), .A2(G105), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT26), .Z(new_n724));
  NAND4_X1  g299(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n719), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n704), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n552), .B2(new_n704), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(new_n730), .B2(G1341), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n714), .A2(new_n718), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n706), .A2(new_n707), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n702), .A2(G2072), .B1(new_n713), .B2(new_n712), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n708), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G4), .A2(G16), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT89), .Z(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n610), .B2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT90), .B(G1348), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n709), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT92), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g318(.A(G140), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT91), .B1(new_n696), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n468), .A2(new_n746), .A3(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n478), .A2(G128), .ZN(new_n748));
  OR2_X1    g323(.A1(G104), .A2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n727), .A2(new_n728), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n709), .B1(new_n758), .B2(G28), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .C1(new_n635), .C2(new_n709), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n717), .A2(G2084), .B1(G1341), .B2(new_n730), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n754), .A2(new_n755), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G21), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G168), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n740), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n704), .A2(G20), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n769), .B(new_n770), .C1(G299), .C2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G164), .A2(new_n709), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G27), .B2(new_n709), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n735), .A2(new_n768), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G303), .A2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(G16), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G1971), .ZN(new_n785));
  INV_X1    g360(.A(G288), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G23), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT33), .B(G1976), .Z(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n782), .B(new_n792), .C1(G16), .C2(new_n783), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n787), .B(new_n789), .C1(G16), .C2(G23), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n785), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n704), .B1(new_n584), .B2(new_n585), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n704), .A2(G6), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n795), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n478), .ZN(new_n805));
  INV_X1    g380(.A(G119), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT86), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT86), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n468), .A2(G131), .ZN(new_n809));
  OR2_X1    g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n802), .B2(new_n803), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n704), .B1(new_n595), .B2(new_n596), .ZN(new_n817));
  INV_X1    g392(.A(G24), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(G16), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT87), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(KEYINPUT87), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n820), .A2(G1986), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(G1986), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT88), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n816), .B(KEYINPUT88), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n804), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g405(.A(KEYINPUT36), .B(new_n804), .C1(new_n826), .C2(new_n827), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n781), .B1(new_n830), .B2(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(G150), .A2(KEYINPUT96), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(new_n781), .C1(new_n830), .C2(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n610), .A2(G559), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n568), .A2(G93), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT97), .B(G55), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(new_n512), .B2(new_n841), .C1(new_n501), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n552), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n839), .A2(new_n844), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n845), .A2(new_n846), .A3(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(G860), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  XNOR2_X1  g426(.A(G164), .B(new_n751), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n701), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n701), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n726), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n726), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n812), .B(new_n627), .ZN(new_n859));
  OR2_X1    g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(G2104), .C1(G118), .C2(new_n477), .ZN(new_n861));
  INV_X1    g436(.A(G142), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n696), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G130), .B2(new_n478), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n851), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n853), .A2(new_n854), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n725), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n868), .B2(new_n855), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT98), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n865), .A3(new_n855), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT99), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n868), .A2(new_n873), .A3(new_n865), .A4(new_n855), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n866), .A2(new_n870), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n635), .B(new_n475), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n483), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n869), .A2(new_n877), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n844), .B(KEYINPUT100), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n623), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n621), .B(KEYINPUT79), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n608), .A2(new_n566), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n602), .B(new_n607), .C1(new_n565), .C2(new_n562), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n566), .A2(new_n608), .A3(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n892), .B2(KEYINPUT101), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(KEYINPUT41), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT102), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n897), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n886), .A2(new_n888), .A3(new_n892), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n883), .B(new_n899), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G290), .A2(new_n786), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(G290), .A2(new_n786), .ZN(new_n907));
  AOI21_X1  g482(.A(G303), .B1(new_n584), .B2(new_n585), .ZN(new_n908));
  NOR2_X1   g483(.A1(G305), .A2(G166), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n907), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n908), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n905), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n903), .B1(new_n900), .B2(new_n901), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n915), .B2(new_n898), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n904), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n904), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n843), .A2(new_n613), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  AND2_X1   g497(.A1(new_n910), .A2(new_n913), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n545), .A2(G651), .A3(new_n570), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(KEYINPUT103), .A3(new_n569), .ZN(new_n925));
  NAND2_X1  g500(.A1(G168), .A2(new_n925), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT103), .B(KEYINPUT104), .C1(new_n924), .C2(new_n569), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(G301), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(G171), .A2(KEYINPUT103), .B1(new_n526), .B2(new_n532), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT104), .B1(G171), .B2(KEYINPUT103), .ZN(new_n933));
  NAND3_X1  g508(.A1(G301), .A2(new_n929), .A3(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n931), .A2(new_n935), .A3(new_n844), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n844), .B1(new_n931), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n897), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n844), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n933), .A2(new_n934), .B1(G168), .B2(new_n925), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n931), .A2(new_n935), .A3(new_n844), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n936), .A2(KEYINPUT105), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n893), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g524(.A(KEYINPUT106), .B(new_n893), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n923), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n944), .A2(new_n943), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n936), .A2(new_n937), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT106), .B1(new_n954), .B2(new_n893), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n947), .A2(new_n948), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n914), .A3(new_n956), .A4(new_n938), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT107), .B1(new_n893), .B2(KEYINPUT41), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n892), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n945), .A2(new_n967), .A3(new_n946), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n953), .A2(new_n892), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n923), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n957), .A2(new_n961), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n957), .A2(new_n971), .A3(new_n974), .A4(new_n961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n960), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n951), .A2(new_n957), .A3(new_n961), .A4(new_n958), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n957), .A2(new_n971), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n980), .B(KEYINPUT44), .C1(new_n961), .C2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(G397));
  OR2_X1    g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n751), .B(new_n753), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n812), .A2(new_n814), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n725), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n812), .A2(new_n814), .ZN(new_n990));
  AND4_X1   g565(.A1(new_n986), .A2(new_n987), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n492), .B2(new_n496), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n470), .A2(G40), .A3(new_n474), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n995), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n497), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT110), .B(G2090), .Z(new_n1004));
  AND4_X1   g579(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n995), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1971), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n995), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1008), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n998), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1012), .B(new_n1013), .C1(new_n1016), .C2(G1971), .ZN(new_n1017));
  NAND3_X1  g592(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT112), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1010), .A2(G8), .A3(new_n1017), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1021), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n580), .A2(new_n583), .A3(G1981), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n580), .B2(new_n583), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n994), .A2(new_n998), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(G8), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n786), .A2(G1976), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n786), .B2(G1976), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1026), .A2(new_n1028), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1015), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT114), .B(new_n998), .C1(new_n994), .C2(KEYINPUT45), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1008), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n766), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1001), .A2(new_n998), .A3(new_n1003), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT115), .B(G2084), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1048), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G286), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT120), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1059), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1052), .A2(new_n766), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT121), .B(new_n1064), .C1(new_n1067), .C2(new_n1048), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1061), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT62), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1052), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(G2078), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1054), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT124), .B(new_n1076), .C1(new_n1077), .C2(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1075), .A2(new_n1080), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G171), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1069), .A2(new_n1087), .A3(new_n1071), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1073), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n777), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1080), .A2(new_n1090), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT125), .B1(new_n1091), .B2(G171), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1083), .A2(new_n1082), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1016), .A2(new_n777), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT124), .B1(new_n1094), .B2(new_n1076), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(G301), .A4(new_n1090), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(new_n1098), .A3(new_n1085), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1054), .A2(new_n773), .ZN(new_n1102));
  INV_X1    g677(.A(new_n565), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n1103), .B2(KEYINPUT118), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(new_n566), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1007), .A2(new_n1008), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT119), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1102), .A2(new_n1106), .A3(new_n1111), .A4(new_n1108), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1105), .ZN(new_n1115));
  INV_X1    g690(.A(new_n610), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1034), .A2(G2067), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1054), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT61), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1007), .A2(new_n988), .A3(new_n1008), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1034), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n619), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n610), .B(new_n1117), .C1(new_n1054), .C2(new_n1118), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1109), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1119), .A2(new_n1133), .A3(new_n610), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1121), .B1(new_n1122), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1091), .A2(G171), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(KEYINPUT54), .C1(G171), .C2(new_n1084), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1101), .A2(new_n1136), .A3(new_n1072), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1047), .B1(new_n1089), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1070), .A2(G8), .A3(G168), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1058), .A2(new_n1143), .A3(G168), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1010), .A2(G8), .A3(new_n1017), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(new_n1021), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1145), .A2(new_n1026), .A3(new_n1046), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1047), .B1(new_n1144), .B2(new_n1142), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1146), .B1(new_n1150), .B2(KEYINPUT117), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1152), .B(new_n1047), .C1(new_n1144), .C2(new_n1142), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1034), .A2(G8), .ZN(new_n1155));
  INV_X1    g730(.A(G1976), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1036), .A2(new_n1156), .A3(new_n786), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1157), .B2(new_n1029), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1026), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1046), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n997), .B1(new_n1140), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT48), .ZN(new_n1163));
  INV_X1    g738(.A(new_n996), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n985), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1164), .B2(new_n991), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n985), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n986), .B2(new_n726), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n996), .A2(new_n988), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT47), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n986), .A2(new_n989), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1175), .A2(new_n987), .B1(G2067), .B2(new_n751), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1168), .B(new_n1174), .C1(new_n996), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n1180));
  NOR2_X1   g754(.A1(G227), .A2(new_n461), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n690), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1180), .B1(G401), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n1184), .A2(KEYINPUT126), .A3(new_n690), .A4(new_n1181), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n878), .B2(new_n880), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n976), .A2(new_n1187), .ZN(G225));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g763(.A1(G225), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n976), .A2(new_n1187), .A3(KEYINPUT127), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1191), .ZN(G308));
endmodule


