//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AOI21_X1  g004(.A(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n188), .A2(new_n190), .A3(G128), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n192), .B2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n189), .B(G146), .C1(new_n193), .C2(new_n194), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n200), .B2(G137), .ZN(new_n205));
  AOI21_X1  g019(.A(G131), .B1(new_n200), .B2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n196), .A2(new_n197), .B1(new_n209), .B2(KEYINPUT68), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n209), .A2(KEYINPUT68), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT2), .B(G113), .Z(new_n212));
  XNOR2_X1  g026(.A(G116), .B(G119), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n212), .A2(KEYINPUT66), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G116), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT2), .B(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(KEYINPUT66), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n188), .A2(new_n190), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  XNOR2_X1  g044(.A(G143), .B(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n226), .ZN(new_n232));
  AND4_X1   g046(.A1(new_n230), .A2(new_n188), .A3(new_n190), .A4(new_n226), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n205), .A2(new_n207), .A3(new_n201), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n208), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(new_n229), .C1(new_n232), .C2(new_n233), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n235), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT28), .B1(new_n224), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n210), .A2(new_n211), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n223), .A2(new_n214), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n247), .A2(new_n248), .B1(new_n241), .B2(new_n224), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n248), .B2(new_n247), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n242), .B1(new_n250), .B2(KEYINPUT28), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(G902), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n189), .A2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n187), .A2(G143), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n195), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n188), .A2(new_n190), .A3(G128), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n197), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT11), .B1(new_n198), .B2(G134), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n272), .A2(new_n206), .B1(new_n236), .B2(G131), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n269), .A2(new_n209), .B1(new_n234), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n246), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n261), .B2(new_n275), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n281), .B2(new_n242), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n282), .A3(new_n256), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT30), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n245), .B1(new_n274), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n261), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n257), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n258), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n293));
  OAI21_X1  g107(.A(G472), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n257), .B1(new_n224), .B2(new_n241), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n287), .A2(new_n297), .A3(new_n300), .A4(new_n296), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n188), .A2(new_n190), .A3(new_n226), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT64), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n231), .A2(new_n230), .A3(new_n226), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n305), .A2(new_n306), .B1(new_n225), .B2(new_n228), .ZN(new_n307));
  INV_X1    g121(.A(G131), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n199), .B2(new_n201), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n272), .B2(new_n206), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n307), .A2(new_n238), .B1(new_n268), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n246), .B1(new_n311), .B2(KEYINPUT30), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n285), .B1(new_n210), .B2(new_n211), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n241), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n261), .A2(new_n256), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(KEYINPUT31), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n256), .B1(new_n279), .B2(new_n282), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT72), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n242), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n278), .B1(new_n277), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n281), .A2(KEYINPUT71), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n257), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n318), .A4(new_n302), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n295), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  AOI211_X1 g145(.A(KEYINPUT32), .B(new_n331), .C1(new_n321), .C2(new_n327), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n294), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT75), .B(G217), .Z(new_n334));
  INV_X1    g148(.A(G902), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(G234), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT80), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(G119), .B(G128), .Z(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n216), .B2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n347), .B(new_n348), .C1(G119), .C2(new_n262), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n345), .B1(G110), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT77), .B(G125), .Z(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT77), .B(G125), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n353), .A4(new_n354), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(KEYINPUT76), .A3(G125), .ZN(new_n361));
  AND3_X1   g175(.A1(KEYINPUT76), .A2(KEYINPUT77), .A3(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(G140), .B1(KEYINPUT77), .B2(G125), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT16), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n360), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n187), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n356), .A2(new_n359), .B1(new_n367), .B2(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G146), .A3(new_n366), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n351), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(G125), .B(G140), .Z(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G146), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n349), .A2(G110), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n343), .A2(new_n344), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n342), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n369), .A2(new_n187), .ZN(new_n382));
  AOI21_X1  g196(.A(G146), .B1(new_n371), .B2(new_n366), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n350), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n379), .A3(new_n341), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n385), .A3(new_n335), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n336), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n381), .A2(new_n385), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n336), .A2(G902), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  OAI21_X1  g210(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G469), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G140), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n337), .A2(G227), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n196), .B2(new_n197), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G104), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G107), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G101), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT81), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(KEYINPUT81), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n406), .A2(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G101), .B1(new_n411), .B2(new_n407), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n265), .B(new_n423), .C1(new_n266), .C2(new_n267), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n419), .A3(new_n420), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n405), .A2(new_n422), .B1(new_n425), .B2(new_n404), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n409), .B1(new_n411), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n410), .A2(G107), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n415), .B2(new_n417), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT82), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(G101), .C1(new_n428), .C2(new_n430), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n434), .A4(new_n419), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(G101), .C1(new_n428), .C2(new_n430), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n235), .A2(new_n240), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n426), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n426), .B(new_n442), .C1(new_n436), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n238), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n238), .B(KEYINPUT83), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n426), .B(new_n445), .C1(new_n436), .C2(new_n439), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n403), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n403), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n269), .A2(new_n421), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n425), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT12), .B1(new_n451), .B2(new_n238), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n453), .B(new_n273), .C1(new_n450), .C2(new_n425), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n399), .B(new_n335), .C1(new_n447), .C2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n399), .A2(new_n335), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n446), .B1(new_n454), .B2(new_n452), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n444), .A2(new_n449), .B1(new_n402), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n460), .B2(G469), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n398), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n337), .A3(G214), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n189), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n252), .B(G214), .C1(KEYINPUT89), .C2(G143), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n308), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n470), .A2(KEYINPUT91), .A3(G131), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT91), .B1(new_n470), .B2(G131), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n463), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(KEYINPUT91), .A3(G131), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(KEYINPUT17), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n370), .A2(new_n473), .A3(new_n476), .A4(new_n372), .ZN(new_n477));
  XNOR2_X1  g291(.A(G113), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(new_n410), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G146), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(G146), .B2(new_n374), .ZN(new_n482));
  AND2_X1   g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n470), .A2(new_n484), .A3(new_n483), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n470), .B2(new_n483), .ZN(new_n486));
  OAI221_X1 g300(.A(new_n482), .B1(new_n470), .B2(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n477), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n479), .B1(new_n477), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n335), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G475), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n480), .A2(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(KEYINPUT19), .B2(new_n374), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n495), .A2(G146), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n372), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  INV_X1    g312(.A(new_n479), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n477), .A2(new_n479), .A3(new_n487), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT20), .B(new_n505), .C1(new_n500), .C2(new_n501), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n491), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G478), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n218), .A2(G122), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT93), .B1(new_n510), .B2(KEYINPUT14), .ZN(new_n511));
  INV_X1    g325(.A(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G116), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(KEYINPUT14), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n510), .A2(KEYINPUT93), .A3(KEYINPUT14), .ZN(new_n516));
  OAI21_X1  g330(.A(G107), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n510), .A3(new_n406), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G134), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n519), .A2(G134), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n262), .A2(G143), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n200), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n513), .A2(new_n510), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G107), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n528), .A2(KEYINPUT92), .A3(new_n518), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT92), .B1(new_n528), .B2(new_n518), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n334), .A2(G953), .A3(new_n396), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n522), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n335), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n537), .B2(new_n335), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n509), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n541), .A2(new_n509), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n507), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n462), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n223), .A2(new_n214), .A3(new_n438), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n434), .A2(KEYINPUT4), .A3(new_n419), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n432), .ZN(new_n551));
  OAI21_X1  g365(.A(G113), .B1(new_n217), .B2(KEYINPUT5), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n213), .A2(KEYINPUT5), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND4_X1   g369(.A1(new_n215), .A2(new_n555), .A3(new_n419), .A4(new_n420), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n548), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n223), .A2(new_n214), .A3(new_n438), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n435), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n547), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n560), .A3(KEYINPUT6), .ZN(new_n561));
  OR3_X1    g375(.A1(new_n559), .A2(KEYINPUT6), .A3(new_n547), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n268), .A2(new_n352), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n229), .B(new_n357), .C1(new_n232), .C2(new_n233), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G224), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT85), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n565), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT7), .B1(new_n566), .B2(G953), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n564), .A3(new_n571), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n559), .B2(new_n547), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n547), .B(KEYINPUT8), .Z(new_n577));
  NOR2_X1   g391(.A1(new_n220), .A2(new_n221), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n554), .B2(new_n553), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n421), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n552), .A2(KEYINPUT86), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n552), .A2(KEYINPUT86), .B1(new_n213), .B2(KEYINPUT5), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n421), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n580), .B(KEYINPUT87), .C1(new_n421), .C2(new_n583), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n576), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G210), .B1(G237), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n570), .A2(new_n589), .A3(new_n591), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT88), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  OAI21_X1  g411(.A(G214), .B1(G237), .B2(G902), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n337), .A2(G952), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT21), .B(G898), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n546), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n333), .A2(new_n395), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT95), .B(G101), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G3));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n321), .B2(new_n327), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(KEYINPUT96), .B(G902), .C1(new_n321), .C2(new_n327), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n328), .A2(new_n335), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT96), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n613), .A2(new_n614), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(KEYINPUT97), .A3(G472), .A4(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT69), .B1(new_n287), .B2(new_n297), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(KEYINPUT31), .B1(new_n299), .B2(new_n301), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n326), .B1(new_n625), .B2(new_n325), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n329), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n462), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n394), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n617), .A2(new_n621), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n538), .A2(G478), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n508), .A2(new_n335), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(G478), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n502), .A2(new_n503), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT20), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n502), .A2(new_n492), .A3(new_n503), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n638), .B1(new_n642), .B2(new_n491), .ZN(new_n643));
  INV_X1    g457(.A(new_n598), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n593), .B2(new_n594), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n606), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n631), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n640), .A2(new_n650), .A3(new_n641), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n506), .A2(KEYINPUT98), .B1(new_n490), .B2(G475), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n544), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n606), .A3(new_n645), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND2_X1  g473(.A1(new_n384), .A2(new_n379), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n392), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n390), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n546), .A2(new_n607), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n617), .A2(new_n621), .A3(new_n628), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NAND2_X1  g483(.A1(new_n664), .A2(new_n645), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n337), .A2(G900), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(G902), .A3(new_n600), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n601), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n670), .A2(new_n654), .A3(new_n653), .A4(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n333), .A2(new_n678), .A3(new_n462), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT100), .B(G128), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G30));
  NAND2_X1  g495(.A1(new_n595), .A2(new_n597), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT38), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n390), .A2(new_n598), .A3(new_n663), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n507), .A2(new_n544), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n595), .A2(new_n687), .A3(new_n597), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n676), .B(KEYINPUT39), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n690), .B1(new_n462), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n462), .A2(new_n690), .A3(new_n691), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n250), .A2(new_n257), .ZN(new_n695));
  INV_X1    g509(.A(new_n624), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n335), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G472), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n330), .B2(new_n332), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n693), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  AND2_X1   g515(.A1(new_n634), .A2(new_n637), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n507), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n677), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n670), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n333), .A2(new_n462), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n628), .A2(KEYINPUT32), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n331), .B1(new_n321), .B2(new_n327), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n295), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n394), .B1(new_n712), .B2(new_n294), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n335), .B1(new_n447), .B2(new_n456), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n397), .A3(new_n457), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n646), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NOR2_X1   g534(.A1(new_n656), .A2(new_n716), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND2_X1  g537(.A1(new_n545), .A2(new_n606), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n716), .A2(new_n724), .A3(new_n670), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n333), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR2_X1   g541(.A1(new_n251), .A2(new_n256), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n329), .B1(new_n728), .B2(new_n319), .ZN(new_n729));
  INV_X1    g543(.A(G472), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n395), .B(new_n729), .C1(new_n613), .C2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n645), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n716), .A2(new_n733), .A3(new_n605), .A4(new_n685), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT101), .B(G122), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G24));
  OAI211_X1 g551(.A(new_n664), .B(new_n729), .C1(new_n613), .C2(new_n730), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n716), .A2(new_n733), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n704), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  AOI21_X1  g556(.A(new_n644), .B1(new_n595), .B2(new_n597), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n462), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n743), .B2(new_n462), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n333), .A3(new_n395), .A4(new_n704), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NOR3_X1   g567(.A1(new_n653), .A2(new_n654), .A3(new_n677), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n747), .A2(new_n333), .A3(new_n395), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND3_X1  g570(.A1(new_n617), .A2(new_n621), .A3(new_n628), .ZN(new_n757));
  INV_X1    g571(.A(new_n507), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n702), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n760), .A2(new_n664), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n757), .A2(KEYINPUT44), .A3(new_n762), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n273), .B1(new_n440), .B2(KEYINPUT84), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n448), .B1(new_n768), .B2(new_n443), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n403), .B1(new_n455), .B2(new_n446), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n444), .A2(new_n449), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n459), .A2(new_n402), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT45), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n774), .A3(G469), .ZN(new_n775));
  INV_X1    g589(.A(new_n458), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT46), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT104), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n457), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n773), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n399), .B1(new_n781), .B2(new_n767), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n458), .B1(new_n782), .B2(new_n774), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n397), .B(new_n691), .C1(new_n780), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n743), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n765), .A2(new_n766), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND3_X1  g604(.A1(new_n704), .A2(new_n743), .A3(new_n394), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n333), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT47), .B(new_n397), .C1(new_n780), .C2(new_n784), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT104), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n795));
  INV_X1    g609(.A(new_n457), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n778), .A2(new_n779), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT47), .B1(new_n799), .B2(new_n397), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n792), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT105), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n397), .B1(new_n780), .B2(new_n784), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n793), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT105), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n792), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n747), .A2(new_n704), .A3(new_n739), .ZN(new_n812));
  INV_X1    g626(.A(new_n743), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n629), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n653), .A2(new_n544), .A3(new_n677), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n333), .A2(new_n664), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n755), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n750), .B2(new_n751), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n333), .A2(new_n725), .B1(new_n732), .B2(new_n734), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n333), .B(new_n395), .C1(new_n721), .C2(new_n717), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n667), .A2(new_n819), .A3(new_n609), .A4(new_n820), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n703), .A2(KEYINPUT108), .B1(new_n507), .B2(new_n654), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n643), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n607), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n631), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n715), .A2(new_n457), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n397), .A3(new_n645), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n738), .A2(new_n831), .A3(new_n705), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n629), .B1(new_n712), .B2(new_n294), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n678), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n733), .A2(new_n664), .A3(new_n685), .A4(new_n677), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n699), .A2(new_n462), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n835), .A3(new_n707), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n679), .A2(new_n707), .A3(new_n837), .A4(new_n741), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n818), .A2(new_n829), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(new_n821), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n615), .A2(new_n616), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n710), .B1(new_n846), .B2(KEYINPUT97), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n617), .A3(new_n630), .A4(new_n826), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n755), .A2(new_n812), .A3(new_n816), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n752), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n679), .A2(new_n707), .A3(new_n741), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n679), .A2(new_n741), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n837), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n838), .A3(new_n840), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n844), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n811), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n853), .A2(new_n838), .A3(new_n840), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n752), .A2(new_n849), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n609), .A2(new_n726), .A3(new_n735), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n859), .A3(new_n667), .A4(new_n820), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n861), .A3(KEYINPUT53), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n841), .A2(new_n842), .ZN(new_n863));
  XNOR2_X1  g677(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n760), .A2(new_n602), .A3(new_n761), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT111), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n682), .A2(new_n870), .A3(new_n598), .A4(new_n732), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n830), .A2(new_n398), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n805), .A2(new_n793), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n683), .A2(new_n688), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n644), .A3(new_n397), .A4(new_n830), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n870), .A2(new_n878), .A3(new_n732), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT50), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT50), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n813), .A2(new_n716), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT116), .Z(new_n887));
  INV_X1    g701(.A(new_n699), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n394), .A2(new_n601), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n758), .A2(new_n638), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n870), .A3(new_n739), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n874), .A2(new_n884), .A3(new_n885), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n870), .A3(new_n713), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT48), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n870), .A2(new_n732), .A3(new_n740), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT117), .Z(new_n899));
  NAND4_X1  g713(.A1(new_n887), .A2(new_n643), .A3(new_n888), .A4(new_n889), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n599), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n895), .A2(new_n897), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n806), .A2(KEYINPUT112), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n806), .A2(KEYINPUT112), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n872), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n871), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT113), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n884), .A2(new_n885), .A3(new_n894), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(KEYINPUT113), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n902), .B1(new_n910), .B2(new_n867), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n866), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(G952), .B2(G953), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n395), .A2(new_n598), .A3(new_n397), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  INV_X1    g729(.A(new_n759), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT49), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(new_n830), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n830), .A2(new_n917), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n875), .A3(new_n888), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n913), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n337), .A2(G952), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n850), .A2(new_n854), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n924), .A2(KEYINPUT53), .B1(new_n841), .B2(new_n842), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT120), .B1(new_n925), .B2(new_n335), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n862), .A2(new_n863), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n928), .A3(G902), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n592), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n561), .A2(new_n562), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n569), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n923), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n335), .B1(new_n862), .B2(new_n863), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(KEYINPUT119), .A3(G210), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT119), .B1(new_n937), .B2(G210), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n936), .A2(new_n942), .ZN(G51));
  INV_X1    g757(.A(new_n775), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n926), .A2(new_n944), .A3(new_n929), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n447), .A2(new_n456), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n458), .B(KEYINPUT121), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT57), .Z(new_n949));
  AOI21_X1  g763(.A(new_n864), .B1(new_n862), .B2(new_n863), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n865), .B2(new_n950), .ZN(new_n951));
  AOI22_X1  g765(.A1(new_n945), .A2(new_n946), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n926), .A2(KEYINPUT122), .A3(new_n944), .A4(new_n929), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n923), .B1(new_n952), .B2(new_n953), .ZN(G54));
  AND2_X1   g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n926), .A2(new_n929), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n500), .A3(new_n501), .ZN(new_n957));
  INV_X1    g771(.A(new_n923), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n926), .A2(new_n502), .A3(new_n929), .A4(new_n955), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n635), .A2(new_n636), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n633), .B(KEYINPUT59), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n864), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n927), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(new_n923), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n963), .B1(new_n856), .B2(new_n865), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n636), .A3(new_n635), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n865), .A2(new_n950), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT123), .B(new_n958), .C1(new_n972), .C2(new_n964), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n925), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n662), .B(KEYINPUT124), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n958), .B1(new_n978), .B2(new_n391), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n978), .A2(new_n391), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n984), .A2(KEYINPUT61), .A3(new_n958), .A4(new_n980), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(G66));
  OAI21_X1  g800(.A(G953), .B1(new_n604), .B2(new_n566), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n829), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n931), .B1(G898), .B2(new_n337), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  OAI21_X1  g804(.A(new_n284), .B1(KEYINPUT30), .B2(new_n311), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(new_n495), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n787), .B1(new_n763), .B2(new_n764), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n766), .A2(new_n993), .B1(new_n802), .B2(new_n808), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n733), .A2(new_n685), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n786), .A2(new_n713), .A3(new_n995), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n752), .A2(new_n755), .A3(new_n851), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n998), .B2(new_n671), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n743), .A2(new_n462), .A3(new_n691), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n825), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(new_n333), .A3(new_n395), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n834), .A2(KEYINPUT62), .A3(new_n700), .A4(new_n707), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n700), .A2(new_n679), .A3(new_n707), .A4(new_n741), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n994), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT126), .B1(new_n1010), .B2(new_n992), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1004), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n809), .A3(new_n789), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n337), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  INV_X1    g830(.A(new_n992), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n999), .A2(new_n1011), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT127), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n999), .A2(new_n1011), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1023), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(G72));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n1014), .B2(new_n860), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1029), .A2(new_n256), .A3(new_n288), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n624), .A2(new_n289), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n1028), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n855), .B2(new_n843), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n994), .A2(new_n997), .A3(new_n829), .ZN(new_n1034));
  AOI211_X1 g848(.A(new_n256), .B(new_n288), .C1(new_n1034), .C2(new_n1028), .ZN(new_n1035));
  NOR4_X1   g849(.A1(new_n1030), .A2(new_n1033), .A3(new_n1035), .A4(new_n923), .ZN(G57));
endmodule


