//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g0011(.A1(G68), .A2(G238), .ZN(new_n212));
  AND2_X1   g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  NOR4_X1   g0013(.A1(new_n208), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n203), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT0), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n231), .A2(new_n233), .A3(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n226), .A2(new_n227), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n228), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT64), .Z(new_n237));
  NOR2_X1   g0037(.A1(new_n224), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n210), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n221), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n209), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n257), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(G77), .C2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n264), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n262), .B(new_n267), .C1(new_n216), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G190), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n230), .B1(new_n232), .B2(new_n215), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT8), .A2(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT8), .A2(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n230), .A2(G33), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n278), .B1(new_n279), .B2(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n229), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n215), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n288), .B1(new_n263), .B2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n289), .A2(KEYINPUT9), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n286), .A2(new_n288), .B1(new_n215), .B2(new_n293), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(KEYINPUT70), .A3(KEYINPUT9), .A4(new_n296), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n275), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n296), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n272), .A2(G200), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n302), .A2(new_n305), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n275), .B(new_n307), .C1(new_n299), .C2(new_n301), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n305), .A4(new_n306), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n272), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n303), .B(new_n316), .C1(G179), .C2(new_n272), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G226), .A2(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n221), .A2(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n256), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n266), .B1(new_n324), .B2(new_n261), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n270), .A2(G238), .A3(new_n264), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n270), .B1(new_n322), .B2(new_n323), .ZN(new_n329));
  NOR4_X1   g0129(.A1(new_n329), .A2(KEYINPUT13), .A3(new_n326), .A4(new_n266), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT14), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n319), .B1(new_n221), .B2(G1698), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n256), .B1(G33), .B2(G97), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n327), .B(new_n267), .C1(new_n270), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n333), .B(KEYINPUT13), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n336), .B2(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n325), .A2(KEYINPUT73), .A3(new_n327), .A4(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(G179), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(G169), .C1(new_n328), .C2(new_n330), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n332), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n295), .ZN(new_n346));
  INV_X1    g0146(.A(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT75), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT75), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n295), .A2(new_n349), .A3(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n291), .A2(G20), .A3(new_n347), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT12), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT76), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n215), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT74), .B1(new_n281), .B2(new_n215), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n230), .C2(G68), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n285), .A2(new_n217), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n288), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT11), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n345), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n338), .A2(new_n339), .A3(G190), .A4(new_n341), .ZN(new_n367));
  OAI21_X1  g0167(.A(G200), .B1(new_n328), .B2(new_n330), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n358), .A2(new_n367), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n282), .A2(new_n280), .A3(new_n283), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G20), .A2(G77), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n285), .C2(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n288), .B1(new_n295), .B2(G77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n293), .A2(new_n217), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT69), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT67), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT68), .B(G107), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G33), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n256), .A2(KEYINPUT67), .A3(G232), .A4(new_n257), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n383), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n261), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n271), .A2(new_n218), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n394), .A2(G190), .A3(new_n267), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n266), .B(new_n395), .C1(new_n393), .C2(new_n261), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n380), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n314), .A2(new_n317), .A3(new_n370), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT79), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT77), .B1(new_n386), .B2(G33), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n259), .A2(new_n257), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n216), .A2(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n387), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n261), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n267), .B1(new_n271), .B2(new_n221), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(G200), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n270), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n416), .A2(G190), .A3(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n402), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n273), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n398), .B1(new_n416), .B2(new_n413), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(KEYINPUT79), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n404), .B1(KEYINPUT3), .B2(new_n268), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n386), .A2(KEYINPUT77), .A3(G33), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n387), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n230), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n403), .B2(new_n405), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT7), .B1(new_n430), .B2(G20), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n431), .A3(G68), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n220), .A2(new_n347), .ZN(new_n433));
  OAI21_X1  g0233(.A(G20), .B1(new_n433), .B2(new_n232), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n280), .A2(G159), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(KEYINPUT16), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n389), .B(new_n230), .C1(KEYINPUT78), .C2(KEYINPUT7), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n256), .B2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n347), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n439), .B1(new_n443), .B2(new_n436), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n438), .A2(new_n288), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n293), .A2(new_n284), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n346), .B2(new_n284), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n423), .A2(new_n449), .A3(KEYINPUT17), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT17), .B1(new_n423), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n445), .A2(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n419), .A2(G179), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n315), .B2(new_n419), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n394), .A2(new_n267), .A3(new_n396), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n315), .ZN(new_n460));
  INV_X1    g0260(.A(new_n379), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n377), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n460), .B(new_n462), .C1(G179), .C2(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n401), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n207), .A2(new_n257), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n430), .B(new_n467), .C1(G264), .C2(new_n257), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n389), .A2(G303), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n261), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n261), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G270), .ZN(new_n476));
  XOR2_X1   g0276(.A(KEYINPUT5), .B(G41), .Z(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(G274), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n471), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n293), .A2(new_n209), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n287), .A2(new_n229), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n263), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n292), .A3(G116), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n209), .A2(G20), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n288), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n230), .C1(G33), .C2(new_n206), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT20), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n288), .A3(new_n486), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n482), .B(new_n485), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n481), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n270), .B1(new_n468), .B2(new_n469), .ZN(new_n497));
  INV_X1    g0297(.A(new_n476), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n497), .A2(new_n498), .A3(new_n479), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT21), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n492), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n483), .A2(new_n292), .A3(new_n484), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(new_n503), .B1(new_n505), .B2(G116), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n315), .B1(new_n506), .B2(new_n482), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n481), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(G190), .ZN(new_n511));
  INV_X1    g0311(.A(new_n494), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n398), .C2(new_n499), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n430), .A2(new_n230), .A3(G68), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n384), .A2(new_n204), .A3(new_n206), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n323), .A2(new_n230), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n285), .A2(KEYINPUT19), .A3(new_n206), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n288), .B1(new_n293), .B2(new_n373), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT84), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n504), .A2(new_n373), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n473), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n270), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n478), .B1(new_n529), .B2(new_n205), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n406), .A2(G238), .A3(new_n257), .A4(new_n387), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n430), .A2(G244), .A3(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n430), .A2(KEYINPUT83), .A3(G238), .A4(new_n257), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n530), .B1(new_n537), .B2(new_n261), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G179), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n315), .B2(new_n538), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n505), .A2(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n522), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n538), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(G200), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(G190), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n527), .A2(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT6), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(new_n550), .B1(new_n206), .B2(G107), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n206), .B2(G107), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n548), .A2(new_n550), .A3(G97), .A4(new_n249), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n440), .A2(new_n442), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n385), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n483), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n504), .A2(new_n206), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n292), .A2(G97), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n387), .A3(new_n388), .A4(G244), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n256), .B2(G250), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n488), .B(new_n565), .C1(new_n566), .C2(new_n257), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT4), .B1(new_n430), .B2(G244), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n387), .A2(new_n388), .A3(G250), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n257), .B1(new_n570), .B2(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n488), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n563), .B1(new_n426), .B2(new_n218), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(KEYINPUT81), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n270), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n479), .B1(new_n475), .B2(G257), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n568), .A2(new_n571), .A3(new_n572), .A4(new_n562), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT81), .B1(new_n573), .B2(new_n574), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n261), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(G190), .A3(new_n577), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n561), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n475), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n480), .B1(new_n586), .B2(new_n207), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n315), .B1(new_n576), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G179), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n577), .B(KEYINPUT82), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n583), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n559), .ZN(new_n592));
  INV_X1    g0392(.A(new_n560), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n554), .A2(G20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n280), .A2(G77), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n594), .A2(new_n557), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n592), .B(new_n593), .C1(new_n596), .C2(new_n483), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n588), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n585), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n230), .A2(KEYINPUT23), .A3(G107), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n204), .A2(G20), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n387), .A3(new_n388), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(KEYINPUT68), .A2(G107), .ZN(new_n606));
  NOR2_X1   g0406(.A1(KEYINPUT68), .A2(G107), .ZN(new_n607));
  OAI21_X1  g0407(.A(G20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT23), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n534), .A2(G20), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n430), .A2(KEYINPUT22), .A3(new_n602), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n600), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n610), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n430), .A2(KEYINPUT22), .A3(new_n602), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(KEYINPUT24), .A3(new_n609), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n288), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n505), .A2(G107), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n292), .A2(G107), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT25), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n406), .A2(G257), .A3(G1698), .A4(new_n387), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G294), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n430), .A2(G250), .A3(new_n257), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n430), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n261), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n479), .B1(new_n475), .B2(G264), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n630), .A2(new_n273), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(G200), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n622), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n315), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n589), .A3(new_n631), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n634), .B2(new_n639), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n546), .B(new_n599), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n466), .A2(new_n514), .A3(new_n643), .ZN(G372));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n543), .A2(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n545), .A3(new_n522), .A4(new_n541), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n585), .A2(new_n647), .A3(new_n634), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n510), .A2(new_n639), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n527), .A2(new_n540), .ZN(new_n651));
  INV_X1    g0451(.A(new_n598), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n645), .A3(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n522), .A2(new_n524), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n540), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n465), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n463), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n369), .A2(new_n660), .B1(new_n345), .B2(new_n365), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n423), .A2(new_n449), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT17), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n423), .A2(new_n449), .A3(KEYINPUT17), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n458), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n314), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n659), .A2(new_n317), .A3(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n291), .A2(new_n230), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n512), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n514), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n510), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n677), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n634), .A2(new_n639), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT86), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n622), .B2(new_n676), .ZN(new_n689));
  INV_X1    g0489(.A(new_n639), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n675), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n679), .A2(new_n676), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n686), .B2(new_n687), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n690), .B2(new_n676), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n225), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G1), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n517), .A2(G116), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n233), .A2(G50), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n702), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n650), .A2(new_n598), .ZN(new_n708));
  INV_X1    g0508(.A(new_n651), .ZN(new_n709));
  OAI221_X1 g0509(.A(new_n657), .B1(new_n645), .B2(new_n647), .C1(new_n655), .C2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT29), .B(new_n676), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n657), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n650), .B2(new_n653), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n675), .B1(new_n713), .B2(new_n655), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n583), .A2(G179), .A3(new_n538), .A4(new_n577), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n630), .A2(new_n471), .A3(new_n476), .A4(new_n631), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n499), .B1(new_n583), .B2(new_n590), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n589), .A3(new_n543), .A4(new_n635), .ZN(new_n722));
  INV_X1    g0522(.A(new_n719), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n576), .A2(new_n587), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n589), .B(new_n530), .C1(new_n537), .C2(new_n261), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n720), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n675), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n514), .A2(new_n675), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n688), .A2(new_n546), .A3(new_n599), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n716), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n707), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n290), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n702), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n684), .B(new_n740), .C1(G330), .C2(new_n681), .ZN(new_n741));
  INV_X1    g0541(.A(new_n681), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n740), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n230), .A2(new_n273), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n589), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n398), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n230), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G58), .A2(new_n750), .B1(new_n754), .B2(G107), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n748), .A2(new_n752), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n747), .A2(new_n751), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n755), .B1(new_n217), .B2(new_n756), .C1(new_n204), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n273), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(G50), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n230), .B1(new_n762), .B2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n206), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n389), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n759), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G68), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n752), .A2(new_n762), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT88), .B(KEYINPUT32), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n761), .A2(new_n765), .A3(new_n767), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n768), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G283), .A2(new_n754), .B1(new_n774), .B2(G329), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT89), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G322), .B2(new_n750), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(G317), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT33), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT33), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n766), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n389), .C1(new_n783), .C2(new_n757), .ZN(new_n784));
  INV_X1    g0584(.A(new_n756), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G311), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n777), .A2(new_n778), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n763), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n773), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n229), .B1(G20), .B2(new_n315), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n256), .A2(G355), .A3(new_n225), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n254), .A2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n430), .A2(new_n700), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G45), .B2(new_n705), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(G116), .B2(new_n225), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n745), .A2(new_n791), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n746), .A2(new_n792), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n741), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  INV_X1    g0602(.A(new_n791), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n430), .B1(new_n804), .B2(new_n768), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n750), .A2(G143), .B1(G150), .B2(new_n766), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  INV_X1    g0607(.A(new_n760), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .C1(new_n769), .C2(new_n756), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  AOI211_X1 g0610(.A(new_n805), .B(new_n810), .C1(G68), .C2(new_n754), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n215), .B2(new_n757), .C1(new_n220), .C2(new_n763), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n749), .A2(new_n788), .B1(new_n768), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n764), .B(new_n814), .C1(G116), .C2(new_n785), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n754), .A2(G87), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n760), .A2(G303), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n389), .B1(new_n757), .B2(new_n249), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G283), .B2(new_n766), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n803), .B1(new_n812), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n803), .A2(new_n744), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT90), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT91), .Z(new_n824));
  AOI211_X1 g0624(.A(new_n740), .B(new_n821), .C1(new_n217), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT92), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n462), .A2(new_n675), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n399), .A2(new_n589), .B1(new_n461), .B2(new_n377), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n400), .A2(new_n827), .B1(new_n828), .B2(new_n460), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(new_n460), .A3(new_n676), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT93), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n380), .A2(new_n397), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n399), .A2(new_n398), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n827), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n463), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT93), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n830), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n826), .B1(new_n744), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n714), .A2(new_n840), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n675), .B(new_n839), .C1(new_n713), .C2(new_n655), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(new_n734), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n740), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT95), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n439), .A2(KEYINPUT94), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n432), .A2(new_n437), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n432), .B2(new_n437), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n850), .A2(new_n851), .A3(new_n483), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n852), .B2(new_n447), .ZN(new_n853));
  INV_X1    g0653(.A(new_n851), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n432), .A2(new_n437), .A3(new_n849), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n288), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(KEYINPUT95), .A3(new_n448), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(new_n455), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n673), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(new_n859), .A3(new_n857), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n860), .A3(new_n662), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  XOR2_X1   g0662(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n453), .B1(new_n455), .B2(new_n859), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n662), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n860), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n456), .A2(new_n457), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT18), .B1(new_n453), .B2(new_n455), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n868), .B1(new_n666), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n866), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n860), .B1(new_n452), .B2(new_n458), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n449), .A2(new_n673), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n666), .B2(new_n871), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n662), .A2(new_n865), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n863), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n866), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT39), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n366), .A2(new_n675), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n365), .A2(new_n675), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n366), .A2(new_n369), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n366), .B2(new_n369), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n658), .A2(new_n676), .A3(new_n840), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n830), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n873), .A2(new_n878), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n898), .A2(new_n899), .B1(new_n871), .B2(new_n673), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT98), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n668), .A2(new_n317), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT99), .B1(new_n715), .B2(new_n466), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT99), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n465), .A4(new_n711), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n904), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n903), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  INV_X1    g0711(.A(new_n887), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n882), .B2(new_n885), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n876), .A2(new_n877), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n727), .A2(new_n675), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT31), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n919));
  INV_X1    g0719(.A(new_n731), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n918), .B(new_n919), .C1(new_n643), .C2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n896), .A2(new_n839), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT40), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n911), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n873), .A2(new_n888), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n832), .B(new_n838), .C1(new_n894), .C2(new_n895), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n730), .B2(new_n732), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n925), .A2(KEYINPUT100), .A3(KEYINPUT40), .A4(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n867), .B2(new_n872), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n876), .A2(new_n877), .A3(new_n874), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n465), .A2(new_n921), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n716), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n910), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n263), .B2(new_n738), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n209), .B1(new_n554), .B2(KEYINPUT35), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n231), .C1(KEYINPUT35), .C2(new_n554), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  OAI21_X1  g0743(.A(G77), .B1(new_n220), .B2(new_n347), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n705), .A2(new_n944), .B1(G50), .B2(new_n347), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(G1), .A3(new_n290), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(new_n943), .A3(new_n946), .ZN(G367));
  INV_X1    g0747(.A(new_n740), .ZN(new_n948));
  INV_X1    g0748(.A(new_n795), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n241), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n798), .B1(new_n225), .B2(new_n373), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n763), .A2(new_n384), .ZN(new_n952));
  INV_X1    g0752(.A(new_n757), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(G116), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT46), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n750), .A2(G303), .B1(G294), .B2(new_n766), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n430), .B1(G97), .B2(new_n754), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G283), .A2(new_n785), .B1(new_n774), .B2(G317), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n952), .B(new_n959), .C1(G311), .C2(new_n760), .ZN(new_n960));
  INV_X1    g0760(.A(new_n763), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(G68), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n279), .B2(new_n749), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n753), .A2(new_n217), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n785), .A2(G50), .B1(G159), .B2(new_n766), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(KEYINPUT108), .ZN(new_n967));
  INV_X1    g0767(.A(G143), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n808), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n389), .B1(new_n953), .B2(G58), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n807), .B2(new_n768), .C1(new_n966), .C2(KEYINPUT108), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n960), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n948), .B1(new_n950), .B2(new_n951), .C1(new_n974), .C2(new_n803), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n542), .A2(new_n675), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n712), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n657), .A2(new_n647), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT101), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n745), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n976), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n739), .A2(G1), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n599), .B1(new_n561), .B2(new_n676), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n652), .A2(new_n675), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT102), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n698), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT44), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(KEYINPUT105), .A3(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n992), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n698), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n991), .A2(KEYINPUT45), .A3(new_n698), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT106), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n694), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1003), .A2(new_n1001), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1008), .A2(new_n995), .A3(new_n1005), .A4(new_n996), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n697), .B1(new_n693), .B2(new_n696), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n684), .B(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1012), .A2(new_n736), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n735), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n987), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n991), .A2(new_n697), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT42), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT43), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n981), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n991), .A2(new_n690), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n675), .B1(new_n1023), .B2(new_n598), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT103), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT103), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n1029), .A3(new_n1022), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n981), .B(KEYINPUT43), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT104), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT104), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n1032), .C1(new_n1019), .C2(new_n1024), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n991), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n695), .A2(new_n1038), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1031), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n985), .B1(new_n1017), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G387));
  NAND2_X1  g0844(.A1(new_n693), .A2(new_n745), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n949), .B1(new_n246), .B2(G45), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n282), .A2(new_n215), .A3(new_n283), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G45), .B1(new_n1047), .B2(KEYINPUT50), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(KEYINPUT50), .B2(new_n1047), .C1(new_n347), .C2(new_n217), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n704), .B(KEYINPUT111), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n704), .A2(new_n225), .A3(new_n256), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G107), .C2(new_n225), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(new_n798), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n953), .A2(G77), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n766), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1055), .B1(new_n215), .B2(new_n749), .C1(new_n1056), .C2(new_n284), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n763), .A2(new_n373), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n785), .A2(G68), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n426), .B1(new_n760), .B2(G159), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G97), .A2(new_n754), .B1(new_n774), .B2(G150), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n749), .A2(new_n779), .B1(new_n756), .B2(new_n783), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT112), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n813), .B2(new_n1056), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G322), .B2(new_n760), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(G283), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n763), .C1(new_n788), .C2(new_n757), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n774), .A2(G326), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n754), .A2(G116), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1073), .A2(new_n426), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1063), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n740), .B(new_n1054), .C1(new_n1078), .C2(new_n791), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1045), .A2(new_n1079), .B1(new_n1012), .B2(new_n986), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n701), .B1(new_n1012), .B2(new_n736), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n1013), .B2(new_n1081), .ZN(G393));
  NAND2_X1  g0882(.A1(new_n251), .A2(new_n795), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1083), .B(new_n798), .C1(new_n206), .C2(new_n225), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n745), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n991), .B2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n756), .A2(new_n284), .B1(new_n768), .B2(new_n968), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n816), .B1(new_n347), .B2(new_n757), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G50), .C2(new_n766), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n808), .A2(new_n279), .B1(new_n749), .B2(new_n769), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n961), .A2(G77), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n430), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1056), .A2(new_n783), .B1(new_n753), .B2(new_n249), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n256), .B(new_n1095), .C1(G116), .C2(new_n961), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n808), .A2(new_n779), .B1(new_n749), .B2(new_n813), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n785), .A2(G294), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n774), .A2(G322), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n757), .A2(new_n1070), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n740), .B(new_n1086), .C1(new_n791), .C2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1010), .B2(new_n986), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n701), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n897), .A2(new_n830), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n896), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n733), .A2(new_n840), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n733), .B2(new_n840), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n676), .B(new_n840), .C1(new_n708), .C2(new_n710), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n830), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1117), .A3(new_n1111), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n465), .A2(G330), .A3(new_n921), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT116), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n909), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n898), .A2(new_n891), .B1(new_n880), .B2(new_n889), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n915), .A2(new_n891), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1117), .B2(new_n896), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1112), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(new_n1111), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1123), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1110), .B1(new_n843), .B2(new_n831), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n891), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n889), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n879), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1116), .A2(new_n830), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n891), .B(new_n915), .C1(new_n1138), .C2(new_n1110), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT115), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n1131), .A3(new_n1111), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1112), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n1122), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1133), .A2(new_n701), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n986), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n890), .A2(new_n744), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n824), .A2(new_n284), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1149), .A2(new_n756), .B1(new_n804), .B2(new_n749), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n389), .B(new_n1150), .C1(G159), .C2(new_n961), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n774), .A2(G125), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n754), .A2(G50), .B1(G128), .B2(new_n760), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n757), .A2(new_n279), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G137), .B2(new_n766), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G87), .A2(new_n953), .B1(new_n785), .B2(G97), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n209), .B2(new_n749), .C1(new_n1070), .C2(new_n808), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n754), .A2(G68), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n774), .A2(G294), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n385), .A2(new_n766), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1093), .A4(new_n1162), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1159), .A2(new_n1163), .A3(new_n256), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT117), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n948), .B(new_n1147), .C1(new_n1166), .C2(new_n803), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1145), .B1(new_n1146), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1144), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n314), .B2(new_n317), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n314), .A2(new_n317), .A3(new_n1173), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n303), .A3(new_n859), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n303), .A2(new_n859), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1176), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n1174), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n934), .A2(new_n924), .A3(new_n928), .A4(G330), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT118), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n929), .A2(KEYINPUT118), .A3(G330), .A4(new_n934), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT119), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT119), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1183), .A2(new_n1181), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n903), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT119), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT119), .ZN(new_n1195));
  AND4_X1   g0995(.A1(new_n903), .A2(new_n1194), .A3(new_n1190), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n909), .A2(new_n1121), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1133), .A2(KEYINPUT121), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT121), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1122), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n1198), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1171), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1194), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n903), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n903), .A2(new_n1194), .A3(new_n1190), .A4(new_n1195), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1203), .A4(new_n1200), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n701), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n986), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT120), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1182), .A2(new_n744), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n426), .B(new_n269), .C1(new_n206), .C2(new_n1056), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n753), .A2(new_n220), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G116), .B2(new_n760), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n962), .A3(new_n1055), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(G107), .C2(new_n750), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n1070), .B2(new_n768), .C1(new_n373), .C2(new_n756), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G41), .B1(new_n774), .B2(G124), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n750), .A2(G128), .B1(new_n961), .B2(G150), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n953), .A2(new_n1148), .B1(G132), .B2(new_n766), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n760), .A2(G125), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n785), .A2(G137), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n268), .B(new_n1223), .C1(new_n1228), .C2(KEYINPUT59), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G159), .B2(new_n754), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n269), .B1(new_n426), .B2(new_n268), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1230), .A2(new_n1231), .B1(new_n215), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n803), .B1(new_n1222), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n823), .A2(G50), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1215), .A2(new_n740), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1213), .A2(new_n1214), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n987), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT120), .B1(new_n1239), .B2(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1212), .A2(new_n1241), .ZN(G375));
  NAND3_X1  g1042(.A1(new_n1198), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1015), .A3(new_n1122), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n740), .B1(new_n824), .B2(new_n347), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1110), .B2(new_n744), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n749), .A2(new_n807), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n808), .A2(new_n804), .B1(new_n757), .B2(new_n769), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n766), .C2(new_n1148), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n774), .A2(G128), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n961), .A2(G50), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n426), .B(new_n1217), .C1(G150), .C2(new_n785), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n757), .A2(new_n206), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n749), .A2(new_n1070), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n965), .B(new_n1255), .C1(new_n385), .C2(new_n785), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n766), .A2(G116), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n256), .B1(new_n774), .B2(G303), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1058), .B1(new_n760), .B2(G294), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1254), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1246), .B1(new_n791), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1119), .B2(new_n986), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1244), .A2(new_n1263), .ZN(G381));
  NOR2_X1   g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT122), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(G390), .A2(G381), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1043), .A3(new_n1267), .A4(new_n1268), .ZN(G407));
  INV_X1    g1069(.A(G213), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1265), .B2(new_n674), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G407), .ZN(G409));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1043), .A2(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1043), .A2(G390), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n801), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT123), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1043), .A2(G390), .A3(new_n1276), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT124), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1043), .A2(G390), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1043), .A2(G390), .A3(new_n1276), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1043), .B2(G390), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1282), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1284), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1212), .A2(new_n1241), .A3(G378), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1197), .A2(new_n1204), .A3(new_n1016), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1213), .A2(new_n1237), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1169), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n701), .B(new_n1122), .C1(new_n1243), .C2(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1243), .A2(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1263), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1270), .A2(G343), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1296), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1296), .A2(new_n1307), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(G2897), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1304), .A2(G2897), .A3(new_n1306), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1308), .A2(KEYINPUT62), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1306), .B(new_n1304), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1291), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1282), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1306), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1323), .B2(new_n1313), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1308), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1273), .B1(new_n1319), .B2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1284), .A2(new_n1290), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1316), .A2(new_n1317), .B1(new_n1323), .B2(new_n1313), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1308), .B2(KEYINPUT62), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1327), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1324), .A2(new_n1308), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1321), .A3(new_n1320), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1333), .A3(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1326), .A2(new_n1334), .ZN(G405));
  NOR2_X1   g1135(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1305), .A2(KEYINPUT127), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1336), .B(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1169), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1292), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G375), .A2(KEYINPUT126), .A3(new_n1169), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1341), .B(new_n1342), .C1(KEYINPUT127), .C2(new_n1305), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1338), .B(new_n1343), .ZN(G402));
endmodule


