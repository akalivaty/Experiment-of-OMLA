

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750;

  XNOR2_X1 U377 ( .A(n455), .B(n454), .ZN(n610) );
  INV_X1 U378 ( .A(G953), .ZN(n734) );
  XNOR2_X1 U379 ( .A(KEYINPUT33), .B(n617), .ZN(n357) );
  NOR2_X2 U380 ( .A1(n733), .A2(n383), .ZN(n375) );
  OR2_X2 U381 ( .A1(n712), .A2(G902), .ZN(n455) );
  NAND2_X2 U382 ( .A1(n413), .A2(n411), .ZN(n733) );
  XNOR2_X2 U383 ( .A(n520), .B(n537), .ZN(n732) );
  XNOR2_X2 U384 ( .A(n478), .B(n431), .ZN(n520) );
  XNOR2_X2 U385 ( .A(n503), .B(KEYINPUT10), .ZN(n532) );
  XNOR2_X2 U386 ( .A(n389), .B(G125), .ZN(n503) );
  NOR2_X1 U387 ( .A1(n546), .A2(n602), .ZN(n514) );
  NOR2_X1 U388 ( .A1(n558), .A2(n650), .ZN(n415) );
  XNOR2_X1 U389 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U390 ( .A(n472), .B(n471), .ZN(n556) );
  XNOR2_X1 U391 ( .A(G101), .B(KEYINPUT66), .ZN(n368) );
  XNOR2_X1 U392 ( .A(n390), .B(KEYINPUT101), .ZN(n374) );
  XNOR2_X1 U393 ( .A(n401), .B(n400), .ZN(n748) );
  XNOR2_X1 U394 ( .A(n561), .B(KEYINPUT19), .ZN(n385) );
  NAND2_X1 U395 ( .A1(n556), .A2(n666), .ZN(n561) );
  BUF_X1 U396 ( .A(n556), .Z(n582) );
  NAND2_X1 U397 ( .A1(n610), .A2(n591), .ZN(n650) );
  XNOR2_X1 U398 ( .A(n416), .B(G469), .ZN(n558) );
  BUF_X1 U399 ( .A(n610), .Z(n399) );
  NOR2_X1 U400 ( .A1(n701), .A2(G902), .ZN(n416) );
  OR2_X1 U401 ( .A1(n628), .A2(G902), .ZN(n425) );
  XNOR2_X1 U402 ( .A(n368), .B(KEYINPUT4), .ZN(n392) );
  XNOR2_X1 U403 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  XNOR2_X1 U404 ( .A(n553), .B(n552), .ZN(n451) );
  AND2_X1 U405 ( .A1(n374), .A2(n744), .ZN(n373) );
  XNOR2_X1 U406 ( .A(n599), .B(KEYINPUT79), .ZN(n600) );
  XNOR2_X1 U407 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U408 ( .A1(n699), .A2(n621), .ZN(n472) );
  XNOR2_X1 U409 ( .A(n657), .B(n424), .ZN(n548) );
  INV_X1 U410 ( .A(KEYINPUT102), .ZN(n424) );
  XNOR2_X1 U411 ( .A(n388), .B(n410), .ZN(n583) );
  INV_X1 U412 ( .A(KEYINPUT39), .ZN(n410) );
  AND2_X1 U413 ( .A1(n516), .A2(n667), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n542), .B(n407), .ZN(n568) );
  XNOR2_X1 U415 ( .A(KEYINPUT13), .B(G475), .ZN(n407) );
  NOR2_X1 U416 ( .A1(n609), .A2(n399), .ZN(n596) );
  XNOR2_X1 U417 ( .A(n512), .B(n358), .ZN(n454) );
  XNOR2_X1 U418 ( .A(n392), .B(n723), .ZN(n477) );
  INV_X1 U419 ( .A(G143), .ZN(n395) );
  XNOR2_X1 U420 ( .A(n732), .B(n430), .ZN(n479) );
  INV_X1 U421 ( .A(G146), .ZN(n430) );
  NAND2_X1 U422 ( .A1(n405), .A2(n357), .ZN(n440) );
  NOR2_X1 U423 ( .A1(n412), .A2(n649), .ZN(n411) );
  INV_X1 U424 ( .A(n743), .ZN(n412) );
  NAND2_X1 U425 ( .A1(n370), .A2(n369), .ZN(n414) );
  XNOR2_X1 U426 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U427 ( .A(n721), .B(n466), .ZN(n467) );
  XNOR2_X1 U428 ( .A(n465), .B(KEYINPUT17), .ZN(n466) );
  INV_X1 U429 ( .A(n558), .ZN(n428) );
  XNOR2_X1 U430 ( .A(n545), .B(n544), .ZN(n684) );
  INV_X1 U431 ( .A(KEYINPUT41), .ZN(n544) );
  XNOR2_X1 U432 ( .A(n486), .B(n485), .ZN(n516) );
  NAND2_X1 U433 ( .A1(n593), .A2(n666), .ZN(n486) );
  XNOR2_X1 U434 ( .A(n387), .B(KEYINPUT22), .ZN(n609) );
  AND2_X1 U435 ( .A1(n592), .A2(n591), .ZN(n404) );
  NAND2_X1 U436 ( .A1(n624), .A2(KEYINPUT72), .ZN(n625) );
  NAND2_X1 U437 ( .A1(n379), .A2(n377), .ZN(n624) );
  NAND2_X1 U438 ( .A1(n710), .A2(G475), .ZN(n436) );
  NAND2_X1 U439 ( .A1(n710), .A2(G210), .ZN(n700) );
  AND2_X1 U440 ( .A1(n670), .A2(n427), .ZN(n426) );
  NAND2_X1 U441 ( .A1(n646), .A2(n564), .ZN(n670) );
  XNOR2_X1 U442 ( .A(KEYINPUT74), .B(G110), .ZN(n418) );
  INV_X1 U443 ( .A(G146), .ZN(n389) );
  XNOR2_X1 U444 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n499) );
  NOR2_X1 U445 ( .A1(G953), .A2(G237), .ZN(n531) );
  XNOR2_X1 U446 ( .A(G137), .B(KEYINPUT5), .ZN(n473) );
  XOR2_X1 U447 ( .A(G113), .B(KEYINPUT93), .Z(n474) );
  XNOR2_X1 U448 ( .A(n445), .B(G104), .ZN(n535) );
  INV_X1 U449 ( .A(G113), .ZN(n445) );
  XOR2_X1 U450 ( .A(KEYINPUT16), .B(G110), .Z(n464) );
  XNOR2_X1 U451 ( .A(n443), .B(G122), .ZN(n521) );
  INV_X1 U452 ( .A(G107), .ZN(n443) );
  XOR2_X1 U453 ( .A(KEYINPUT68), .B(G131), .Z(n537) );
  XNOR2_X1 U454 ( .A(G122), .B(KEYINPUT12), .ZN(n529) );
  XOR2_X1 U455 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n530) );
  XNOR2_X1 U456 ( .A(n419), .B(n417), .ZN(n496) );
  XNOR2_X1 U457 ( .A(n493), .B(n418), .ZN(n417) );
  XNOR2_X1 U458 ( .A(n504), .B(n494), .ZN(n419) );
  XNOR2_X1 U459 ( .A(G104), .B(G107), .ZN(n493) );
  OR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n483) );
  XNOR2_X1 U461 ( .A(n481), .B(G472), .ZN(n482) );
  XNOR2_X1 U462 ( .A(n432), .B(KEYINPUT0), .ZN(n601) );
  NAND2_X1 U463 ( .A1(n385), .A2(n590), .ZN(n432) );
  INV_X1 U464 ( .A(KEYINPUT3), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n444), .B(n441), .ZN(n721) );
  XNOR2_X1 U466 ( .A(n521), .B(n442), .ZN(n441) );
  XNOR2_X1 U467 ( .A(n464), .B(n535), .ZN(n444) );
  INV_X1 U468 ( .A(KEYINPUT70), .ZN(n442) );
  XNOR2_X1 U469 ( .A(n505), .B(n398), .ZN(n397) );
  INV_X1 U470 ( .A(KEYINPUT23), .ZN(n398) );
  XNOR2_X1 U471 ( .A(n532), .B(n504), .ZN(n729) );
  AND2_X1 U472 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U473 ( .A1(n718), .A2(n383), .ZN(n381) );
  INV_X1 U474 ( .A(G134), .ZN(n431) );
  XNOR2_X1 U475 ( .A(n437), .B(KEYINPUT35), .ZN(n619) );
  XNOR2_X1 U476 ( .A(n440), .B(n439), .ZN(n438) );
  INV_X1 U477 ( .A(KEYINPUT34), .ZN(n439) );
  NAND2_X1 U478 ( .A1(n710), .A2(G472), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n510), .B(n509), .ZN(n712) );
  XNOR2_X1 U480 ( .A(n508), .B(n457), .ZN(n509) );
  XNOR2_X1 U481 ( .A(n729), .B(KEYINPUT87), .ZN(n510) );
  XNOR2_X1 U482 ( .A(n397), .B(n506), .ZN(n508) );
  NAND2_X1 U483 ( .A1(n710), .A2(G469), .ZN(n448) );
  AND2_X1 U484 ( .A1(n429), .A2(n428), .ZN(n562) );
  INV_X1 U485 ( .A(KEYINPUT40), .ZN(n400) );
  NOR2_X2 U486 ( .A1(n583), .A2(n564), .ZN(n401) );
  XNOR2_X1 U487 ( .A(n560), .B(KEYINPUT108), .ZN(n745) );
  NOR2_X1 U488 ( .A1(n577), .A2(n561), .ZN(n557) );
  AND2_X1 U489 ( .A1(n596), .A2(n391), .ZN(n598) );
  AND2_X1 U490 ( .A1(n595), .A2(n611), .ZN(n391) );
  AND2_X1 U491 ( .A1(n515), .A2(n396), .ZN(n569) );
  AND2_X1 U492 ( .A1(n516), .A2(n360), .ZN(n396) );
  AND2_X1 U493 ( .A1(n429), .A2(n427), .ZN(n642) );
  OR2_X2 U494 ( .A1(n609), .A2(n386), .ZN(n613) );
  NAND2_X1 U495 ( .A1(n612), .A2(n595), .ZN(n386) );
  XNOR2_X1 U496 ( .A(n706), .B(n408), .ZN(n709) );
  XNOR2_X1 U497 ( .A(n708), .B(n707), .ZN(n408) );
  INV_X1 U498 ( .A(KEYINPUT60), .ZN(n433) );
  INV_X1 U499 ( .A(KEYINPUT56), .ZN(n393) );
  XNOR2_X1 U500 ( .A(KEYINPUT25), .B(KEYINPUT89), .ZN(n358) );
  XOR2_X1 U501 ( .A(n474), .B(n473), .Z(n359) );
  AND2_X1 U502 ( .A1(n568), .A2(n567), .ZN(n360) );
  AND2_X1 U503 ( .A1(n619), .A2(n620), .ZN(n361) );
  BUF_X1 U504 ( .A(n601), .Z(n618) );
  XOR2_X1 U505 ( .A(n628), .B(n627), .Z(n362) );
  XOR2_X1 U506 ( .A(n705), .B(n704), .Z(n363) );
  XOR2_X1 U507 ( .A(n699), .B(n698), .Z(n364) );
  XNOR2_X1 U508 ( .A(n703), .B(n702), .ZN(n365) );
  NOR2_X1 U509 ( .A1(G952), .A2(n734), .ZN(n714) );
  INV_X1 U510 ( .A(n714), .ZN(n421) );
  XOR2_X1 U511 ( .A(n630), .B(n629), .Z(n366) );
  XOR2_X1 U512 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n367) );
  INV_X1 U513 ( .A(n392), .ZN(n495) );
  NAND2_X1 U514 ( .A1(n374), .A2(n361), .ZN(n369) );
  NAND2_X1 U515 ( .A1(n373), .A2(n371), .ZN(n370) );
  XNOR2_X1 U516 ( .A(n372), .B(n600), .ZN(n371) );
  NAND2_X1 U517 ( .A1(n747), .A2(n636), .ZN(n372) );
  INV_X1 U518 ( .A(n619), .ZN(n744) );
  INV_X1 U519 ( .A(n718), .ZN(n382) );
  NAND2_X1 U520 ( .A1(n382), .A2(n375), .ZN(n689) );
  NAND2_X1 U521 ( .A1(n382), .A2(n376), .ZN(n384) );
  INV_X1 U522 ( .A(n733), .ZN(n376) );
  NAND2_X1 U523 ( .A1(n382), .A2(n378), .ZN(n377) );
  NOR2_X1 U524 ( .A1(n733), .A2(n383), .ZN(n378) );
  NAND2_X1 U525 ( .A1(n733), .A2(n383), .ZN(n380) );
  AND2_X1 U526 ( .A1(n384), .A2(n367), .ZN(n691) );
  INV_X1 U527 ( .A(KEYINPUT2), .ZN(n383) );
  AND2_X1 U528 ( .A1(n428), .A2(n385), .ZN(n427) );
  NAND2_X1 U529 ( .A1(n405), .A2(n404), .ZN(n387) );
  XNOR2_X1 U530 ( .A(n423), .B(n362), .ZN(n422) );
  XNOR2_X1 U531 ( .A(n436), .B(n363), .ZN(n435) );
  XNOR2_X1 U532 ( .A(n448), .B(n365), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n415), .B(KEYINPUT91), .ZN(n602) );
  AND2_X4 U534 ( .A1(n626), .A2(n625), .ZN(n710) );
  NAND2_X1 U535 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U536 ( .A1(n435), .A2(n421), .ZN(n434) );
  NAND2_X1 U537 ( .A1(n447), .A2(n421), .ZN(n446) );
  XNOR2_X1 U538 ( .A(n434), .B(n433), .ZN(G60) );
  NAND2_X1 U539 ( .A1(n409), .A2(n515), .ZN(n388) );
  NAND2_X1 U540 ( .A1(n750), .A2(n614), .ZN(n390) );
  XNOR2_X2 U541 ( .A(n613), .B(KEYINPUT100), .ZN(n750) );
  XNOR2_X2 U542 ( .A(n403), .B(n402), .ZN(n723) );
  INV_X1 U543 ( .A(n601), .ZN(n405) );
  XNOR2_X1 U544 ( .A(n477), .B(n478), .ZN(n461) );
  XNOR2_X1 U545 ( .A(n394), .B(n393), .ZN(G51) );
  NAND2_X1 U546 ( .A1(n406), .A2(n421), .ZN(n394) );
  XNOR2_X2 U547 ( .A(n395), .B(G128), .ZN(n478) );
  NOR2_X1 U548 ( .A1(n576), .A2(n453), .ZN(n452) );
  XNOR2_X1 U549 ( .A(n572), .B(n571), .ZN(n573) );
  NOR2_X1 U550 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X2 U551 ( .A(G119), .B(G116), .ZN(n403) );
  INV_X1 U552 ( .A(n479), .ZN(n498) );
  XNOR2_X1 U553 ( .A(n700), .B(n364), .ZN(n406) );
  NAND2_X1 U554 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n541), .B(n540), .ZN(n705) );
  XNOR2_X1 U556 ( .A(n450), .B(n449), .ZN(n413) );
  XNOR2_X2 U557 ( .A(n414), .B(KEYINPUT45), .ZN(n718) );
  XNOR2_X1 U558 ( .A(n420), .B(n366), .ZN(G57) );
  INV_X1 U559 ( .A(n657), .ZN(n604) );
  XNOR2_X2 U560 ( .A(n425), .B(n482), .ZN(n657) );
  XNOR2_X1 U561 ( .A(n549), .B(KEYINPUT28), .ZN(n429) );
  NAND2_X1 U562 ( .A1(n429), .A2(n426), .ZN(n566) );
  NAND2_X1 U563 ( .A1(n438), .A2(n360), .ZN(n437) );
  XNOR2_X1 U564 ( .A(n575), .B(KEYINPUT71), .ZN(n576) );
  XNOR2_X1 U565 ( .A(n446), .B(KEYINPUT119), .ZN(G54) );
  INV_X1 U566 ( .A(KEYINPUT48), .ZN(n449) );
  INV_X1 U567 ( .A(n745), .ZN(n453) );
  AND2_X1 U568 ( .A1(G214), .A2(n531), .ZN(n456) );
  AND2_X1 U569 ( .A1(n522), .A2(G221), .ZN(n457) );
  INV_X1 U570 ( .A(KEYINPUT77), .ZN(n571) );
  XNOR2_X1 U571 ( .A(n495), .B(n496), .ZN(n497) );
  XNOR2_X1 U572 ( .A(n359), .B(n475), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n532), .B(n456), .ZN(n533) );
  XNOR2_X1 U574 ( .A(n498), .B(n497), .ZN(n701) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n480) );
  INV_X1 U576 ( .A(n621), .ZN(n622) );
  INV_X1 U577 ( .A(KEYINPUT73), .ZN(n513) );
  INV_X1 U578 ( .A(KEYINPUT82), .ZN(n629) );
  INV_X1 U579 ( .A(n461), .ZN(n459) );
  AND2_X1 U580 ( .A1(G224), .A2(n734), .ZN(n460) );
  INV_X1 U581 ( .A(n460), .ZN(n458) );
  NAND2_X1 U582 ( .A1(n459), .A2(n458), .ZN(n463) );
  NAND2_X1 U583 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U584 ( .A1(n463), .A2(n462), .ZN(n468) );
  XOR2_X1 U585 ( .A(n503), .B(KEYINPUT18), .Z(n465) );
  XNOR2_X2 U586 ( .A(n468), .B(n467), .ZN(n699) );
  XOR2_X1 U587 ( .A(KEYINPUT83), .B(KEYINPUT75), .Z(n470) );
  NAND2_X1 U588 ( .A1(G210), .A2(n483), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n582), .B(KEYINPUT38), .ZN(n543) );
  NAND2_X1 U590 ( .A1(G210), .A2(n531), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n480), .B(n479), .ZN(n628) );
  INV_X1 U592 ( .A(KEYINPUT69), .ZN(n481) );
  INV_X1 U593 ( .A(n548), .ZN(n593) );
  NAND2_X1 U594 ( .A1(G214), .A2(n483), .ZN(n666) );
  XNOR2_X1 U595 ( .A(KEYINPUT106), .B(KEYINPUT30), .ZN(n484) );
  XNOR2_X1 U596 ( .A(n484), .B(KEYINPUT105), .ZN(n485) );
  NAND2_X1 U597 ( .A1(G234), .A2(G237), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n487), .B(KEYINPUT14), .ZN(n489) );
  NAND2_X1 U599 ( .A1(G952), .A2(n489), .ZN(n682) );
  NOR2_X1 U600 ( .A1(n682), .A2(G953), .ZN(n488) );
  XNOR2_X1 U601 ( .A(n488), .B(KEYINPUT84), .ZN(n587) );
  NAND2_X1 U602 ( .A1(n489), .A2(G902), .ZN(n490) );
  XNOR2_X1 U603 ( .A(n490), .B(KEYINPUT85), .ZN(n585) );
  NAND2_X1 U604 ( .A1(n585), .A2(G953), .ZN(n491) );
  NOR2_X1 U605 ( .A1(G900), .A2(n491), .ZN(n492) );
  NOR2_X1 U606 ( .A1(n587), .A2(n492), .ZN(n546) );
  XOR2_X1 U607 ( .A(G137), .B(G140), .Z(n504) );
  NAND2_X1 U608 ( .A1(G227), .A2(n734), .ZN(n494) );
  NAND2_X1 U609 ( .A1(n621), .A2(G234), .ZN(n500) );
  XNOR2_X1 U610 ( .A(n500), .B(n499), .ZN(n511) );
  NAND2_X1 U611 ( .A1(n511), .A2(G221), .ZN(n501) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(n501), .Z(n502) );
  XNOR2_X1 U613 ( .A(KEYINPUT90), .B(n502), .ZN(n591) );
  XOR2_X1 U614 ( .A(KEYINPUT24), .B(G110), .Z(n506) );
  XNOR2_X1 U615 ( .A(G128), .B(G119), .ZN(n505) );
  NAND2_X1 U616 ( .A1(G234), .A2(n734), .ZN(n507) );
  XOR2_X1 U617 ( .A(KEYINPUT8), .B(n507), .Z(n522) );
  NAND2_X1 U618 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U619 ( .A(KEYINPUT99), .B(G478), .ZN(n528) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n518) );
  XNOR2_X1 U621 ( .A(G116), .B(KEYINPUT7), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U623 ( .A(n520), .B(n519), .ZN(n526) );
  XOR2_X1 U624 ( .A(n521), .B(KEYINPUT98), .Z(n524) );
  NAND2_X1 U625 ( .A1(G217), .A2(n522), .ZN(n523) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n708) );
  NOR2_X1 U628 ( .A1(G902), .A2(n708), .ZN(n527) );
  XNOR2_X1 U629 ( .A(n528), .B(n527), .ZN(n567) );
  INV_X1 U630 ( .A(n567), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n530), .B(n529), .ZN(n534) );
  XOR2_X1 U632 ( .A(n534), .B(n533), .Z(n541) );
  XNOR2_X1 U633 ( .A(G143), .B(n535), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n536), .B(G140), .ZN(n539) );
  XNOR2_X1 U635 ( .A(n537), .B(KEYINPUT95), .ZN(n538) );
  NOR2_X1 U636 ( .A1(G902), .A2(n705), .ZN(n542) );
  NAND2_X1 U637 ( .A1(n563), .A2(n568), .ZN(n564) );
  XOR2_X1 U638 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n551) );
  NOR2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n592) );
  INV_X1 U640 ( .A(n592), .ZN(n669) );
  INV_X1 U641 ( .A(n543), .ZN(n667) );
  NAND2_X1 U642 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U643 ( .A1(n669), .A2(n671), .ZN(n545) );
  NOR2_X1 U644 ( .A1(n546), .A2(n399), .ZN(n547) );
  NAND2_X1 U645 ( .A1(n591), .A2(n547), .ZN(n554) );
  NOR2_X1 U646 ( .A1(n548), .A2(n554), .ZN(n549) );
  NAND2_X1 U647 ( .A1(n684), .A2(n562), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n551), .B(n550), .ZN(n749) );
  NAND2_X1 U649 ( .A1(n748), .A2(n749), .ZN(n553) );
  XOR2_X1 U650 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n552) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(n604), .Z(n595) );
  INV_X1 U652 ( .A(n595), .ZN(n615) );
  XNOR2_X1 U653 ( .A(n564), .B(KEYINPUT103), .ZN(n641) );
  INV_X1 U654 ( .A(n641), .ZN(n644) );
  NOR2_X1 U655 ( .A1(n554), .A2(n644), .ZN(n555) );
  NAND2_X1 U656 ( .A1(n615), .A2(n555), .ZN(n577) );
  XNOR2_X1 U657 ( .A(KEYINPUT36), .B(n557), .ZN(n559) );
  XNOR2_X1 U658 ( .A(n558), .B(KEYINPUT1), .ZN(n651) );
  INV_X1 U659 ( .A(n651), .ZN(n611) );
  NAND2_X1 U660 ( .A1(n559), .A2(n611), .ZN(n560) );
  NOR2_X1 U661 ( .A1(n563), .A2(n568), .ZN(n637) );
  INV_X1 U662 ( .A(n637), .ZN(n646) );
  XOR2_X1 U663 ( .A(KEYINPUT47), .B(KEYINPUT67), .Z(n565) );
  NOR2_X1 U664 ( .A1(n566), .A2(n565), .ZN(n574) );
  NAND2_X1 U665 ( .A1(KEYINPUT47), .A2(n566), .ZN(n570) );
  NAND2_X1 U666 ( .A1(n582), .A2(n569), .ZN(n640) );
  NAND2_X1 U667 ( .A1(n570), .A2(n640), .ZN(n572) );
  XOR2_X1 U668 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n580) );
  NOR2_X1 U669 ( .A1(n611), .A2(n577), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n578), .A2(n666), .ZN(n579) );
  XNOR2_X1 U671 ( .A(n580), .B(n579), .ZN(n581) );
  NOR2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n649) );
  NOR2_X1 U673 ( .A1(n646), .A2(n583), .ZN(n584) );
  XNOR2_X1 U674 ( .A(n584), .B(KEYINPUT109), .ZN(n743) );
  NOR2_X1 U675 ( .A1(G898), .A2(n734), .ZN(n725) );
  NAND2_X1 U676 ( .A1(n585), .A2(n725), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT86), .B(n586), .ZN(n589) );
  INV_X1 U678 ( .A(n587), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U680 ( .A(n591), .ZN(n653) );
  NOR2_X1 U681 ( .A1(n593), .A2(n611), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n596), .A2(n594), .ZN(n636) );
  XNOR2_X1 U683 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n597) );
  XNOR2_X1 U684 ( .A(n598), .B(n597), .ZN(n747) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n620), .A2(KEYINPUT78), .ZN(n599) );
  NOR2_X1 U687 ( .A1(n618), .A2(n602), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n603), .B(KEYINPUT92), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n632) );
  NOR2_X1 U690 ( .A1(n651), .A2(n650), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n657), .A2(n616), .ZN(n662) );
  NOR2_X1 U692 ( .A1(n618), .A2(n662), .ZN(n607) );
  XNOR2_X1 U693 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n606) );
  XNOR2_X1 U694 ( .A(n607), .B(n606), .ZN(n647) );
  NAND2_X1 U695 ( .A1(n632), .A2(n647), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n608), .A2(n670), .ZN(n614) );
  INV_X1 U697 ( .A(n399), .ZN(n654) );
  NOR2_X1 U698 ( .A1(n611), .A2(n654), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n617) );
  INV_X1 U700 ( .A(KEYINPUT72), .ZN(n688) );
  NAND2_X1 U701 ( .A1(n689), .A2(n688), .ZN(n623) );
  AND2_X2 U702 ( .A1(n623), .A2(n622), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT62), .B(KEYINPUT81), .Z(n627) );
  XNOR2_X1 U704 ( .A(KEYINPUT63), .B(KEYINPUT110), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n644), .A2(n632), .ZN(n631) );
  XOR2_X1 U706 ( .A(G104), .B(n631), .Z(G6) );
  NOR2_X1 U707 ( .A1(n646), .A2(n632), .ZN(n634) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U710 ( .A(G107), .B(n635), .ZN(G9) );
  XNOR2_X1 U711 ( .A(G110), .B(n636), .ZN(G12) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U713 ( .A1(n642), .A2(n637), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n639), .B(n638), .ZN(G30) );
  XNOR2_X1 U715 ( .A(G143), .B(n640), .ZN(G45) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(G146), .ZN(G48) );
  NOR2_X1 U718 ( .A1(n647), .A2(n644), .ZN(n645) );
  XOR2_X1 U719 ( .A(G113), .B(n645), .Z(G15) );
  NOR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U721 ( .A(G116), .B(n648), .Z(G18) );
  XOR2_X1 U722 ( .A(G140), .B(n649), .Z(G42) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U724 ( .A(KEYINPUT50), .B(n652), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n656) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n664) );
  XOR2_X1 U731 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U733 ( .A1(n665), .A2(n684), .ZN(n678) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n674) );
  INV_X1 U736 ( .A(n670), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(KEYINPUT113), .B(n675), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n357), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U742 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT52), .B(n680), .Z(n681) );
  NOR2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n683), .B(KEYINPUT115), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n357), .A2(n684), .ZN(n685) );
  NAND2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U748 ( .A(n687), .B(KEYINPUT116), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n734), .A2(n694), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT53), .B(n695), .Z(G75) );
  XOR2_X1 U754 ( .A(KEYINPUT55), .B(KEYINPUT80), .Z(n697) );
  XNOR2_X1 U755 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U757 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT57), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n704) );
  XOR2_X1 U760 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n707) );
  NAND2_X1 U761 ( .A1(n710), .A2(G478), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n714), .A2(n709), .ZN(G63) );
  NAND2_X1 U763 ( .A1(G217), .A2(n710), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(G898), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n717), .B(KEYINPUT123), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n718), .A2(G953), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n727) );
  XOR2_X1 U772 ( .A(G101), .B(n721), .Z(n722) );
  XNOR2_X1 U773 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U775 ( .A(n727), .B(n726), .Z(n728) );
  XNOR2_X1 U776 ( .A(KEYINPUT124), .B(n728), .ZN(G69) );
  XOR2_X1 U777 ( .A(n729), .B(KEYINPUT4), .Z(n730) );
  XNOR2_X1 U778 ( .A(KEYINPUT125), .B(n730), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n732), .B(n731), .ZN(n737) );
  XNOR2_X1 U780 ( .A(n737), .B(n733), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n736), .ZN(n742) );
  XNOR2_X1 U783 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U785 ( .A1(G953), .A2(n739), .ZN(n740) );
  XOR2_X1 U786 ( .A(KEYINPUT127), .B(n740), .Z(n741) );
  NAND2_X1 U787 ( .A1(n742), .A2(n741), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G134), .B(n743), .ZN(G36) );
  XNOR2_X1 U789 ( .A(G122), .B(n744), .ZN(G24) );
  XOR2_X1 U790 ( .A(n745), .B(G125), .Z(n746) );
  XNOR2_X1 U791 ( .A(KEYINPUT37), .B(n746), .ZN(G27) );
  XNOR2_X1 U792 ( .A(G119), .B(n747), .ZN(G21) );
  XNOR2_X1 U793 ( .A(n748), .B(G131), .ZN(G33) );
  XNOR2_X1 U794 ( .A(G137), .B(n749), .ZN(G39) );
  XNOR2_X1 U795 ( .A(n750), .B(G101), .ZN(G3) );
endmodule

