//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT1), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n209), .B(new_n213), .C1(new_n207), .C2(new_n210), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT26), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n218), .A2(new_n224), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT27), .B1(new_n226), .B2(KEYINPUT66), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT67), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT28), .A4(new_n231), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n240), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n231), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n232), .B2(new_n233), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n225), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n217), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n224), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n245), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n249), .B1(new_n257), .B2(KEYINPUT24), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n259));
  OAI221_X1 g058(.A(new_n246), .B1(G183gat), .B2(G190gat), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n224), .A4(new_n254), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n244), .A2(new_n262), .A3(KEYINPUT70), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT70), .B1(new_n244), .B2(new_n262), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n216), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n262), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n215), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n202), .B1(new_n271), .B2(KEYINPUT73), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT34), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n272), .A2(new_n273), .B1(new_n202), .B2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n266), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n244), .A2(new_n262), .A3(KEYINPUT70), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n215), .B1(new_n269), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n264), .A2(new_n216), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n279), .B1(new_n284), .B2(KEYINPUT32), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n266), .B1(new_n265), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n286), .B2(KEYINPUT33), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n284), .B(KEYINPUT32), .C1(new_n289), .C2(new_n279), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n276), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n293), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n298), .B(new_n299), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(KEYINPUT83), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(G141gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n301), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(KEYINPUT84), .A3(new_n301), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n298), .A2(new_n299), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n298), .B2(new_n305), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI211_X1 g121(.A(KEYINPUT85), .B(KEYINPUT2), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n318), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n308), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n312), .A2(KEYINPUT84), .A3(new_n301), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT84), .B1(new_n312), .B2(new_n301), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n308), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n307), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT87), .B1(new_n330), .B2(KEYINPUT3), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT86), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n306), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT29), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G211gat), .B(G218gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT76), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  AND2_X1   g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n343), .A2(KEYINPUT22), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n340), .A2(new_n346), .ZN(new_n349));
  OR3_X1    g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT77), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n334), .B1(new_n356), .B2(new_n336), .ZN(new_n357));
  OAI211_X1 g156(.A(G228gat), .B(G233gat), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n348), .B2(new_n349), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n360), .A2(new_n336), .ZN(new_n361));
  OAI221_X1 g160(.A(new_n359), .B1(new_n334), .B2(new_n361), .C1(new_n338), .C2(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(G22gat), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(G22gat), .B1(new_n358), .B2(new_n362), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT92), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  OAI22_X1  g168(.A1(new_n364), .A2(new_n365), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n365), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n369), .B(KEYINPUT92), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n373), .A3(new_n363), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n297), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT81), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT82), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n267), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n244), .A2(new_n262), .A3(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n267), .A2(new_n355), .A3(new_n386), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n352), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n355), .A3(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n394), .A3(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n267), .A2(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n390), .B1(new_n397), .B2(new_n352), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n392), .A2(KEYINPUT79), .B1(new_n267), .B2(new_n387), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n353), .B1(new_n401), .B2(new_n395), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT80), .B1(new_n402), .B2(new_n390), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n352), .ZN(new_n405));
  INV_X1    g204(.A(new_n381), .ZN(new_n406));
  INV_X1    g205(.A(new_n390), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT30), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n398), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n381), .A2(new_n404), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G1gat), .B(G29gat), .Z(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n216), .B1(new_n334), .B2(new_n336), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n331), .B2(new_n337), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n307), .B(new_n215), .C1(new_n325), .C2(new_n329), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n330), .A2(new_n216), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n420), .ZN(new_n430));
  INV_X1    g229(.A(new_n423), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(KEYINPUT88), .C1(new_n419), .C2(new_n425), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n215), .B1(new_n330), .B2(KEYINPUT3), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n333), .A2(new_n328), .ZN(new_n437));
  AND4_X1   g236(.A1(new_n335), .A2(new_n437), .A3(new_n336), .A4(new_n307), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT88), .B1(new_n441), .B2(new_n432), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n428), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT90), .B(KEYINPUT6), .Z(new_n444));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n431), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n426), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n448), .A2(new_n433), .B1(new_n427), .B2(new_n426), .ZN(new_n449));
  INV_X1    g248(.A(new_n417), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n443), .B(new_n444), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n427), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n434), .B2(new_n442), .ZN(new_n453));
  INV_X1    g252(.A(new_n444), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n417), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n412), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n376), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n417), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n448), .A2(new_n433), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n454), .B1(new_n462), .B2(new_n428), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n460), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n455), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT72), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n291), .A2(new_n292), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n469), .A3(new_n276), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n293), .A2(KEYINPUT72), .B1(new_n274), .B2(new_n275), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT75), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n276), .A2(new_n293), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n370), .B2(new_n374), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n466), .A2(new_n475), .A3(new_n412), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n459), .B1(new_n478), .B2(KEYINPUT35), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n470), .A2(new_n471), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT75), .B1(new_n473), .B2(new_n469), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n296), .A2(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n375), .ZN(new_n488));
  INV_X1    g287(.A(new_n455), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n443), .A2(new_n444), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n450), .B1(new_n462), .B2(new_n452), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT91), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n460), .A2(new_n463), .A3(new_n461), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n404), .A2(new_n381), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n409), .A2(new_n411), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n488), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n430), .B2(new_n431), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n429), .A2(KEYINPUT93), .A3(new_n423), .A4(new_n420), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n422), .A2(new_n424), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n423), .B1(new_n505), .B2(new_n440), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n431), .C1(new_n419), .C2(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n450), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT94), .B(new_n499), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n507), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(KEYINPUT94), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n453), .A2(new_n417), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR4_X1   g313(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n381), .A4(new_n390), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n410), .B1(new_n398), .B2(new_n406), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n406), .B1(new_n400), .B2(new_n403), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n511), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT38), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n404), .A2(KEYINPUT37), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n406), .B1(new_n398), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n397), .A2(new_n353), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n388), .A2(new_n389), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n526), .B2(new_n352), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT38), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n451), .A2(new_n529), .A3(new_n455), .A4(new_n408), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n519), .B(new_n375), .C1(new_n524), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n487), .A2(new_n498), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n480), .A2(KEYINPUT96), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n479), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  AND2_X1   g337(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n546));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(G1gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n558), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n550), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n549), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT18), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(KEYINPUT18), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n562), .B(new_n549), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n564), .B(KEYINPUT13), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT97), .B(KEYINPUT11), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT12), .Z(new_n577));
  OR2_X1    g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(G64gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n582), .A2(G57gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(G57gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n586));
  AND2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n581), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n585), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n562), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n598), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n550), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  INV_X1    g414(.A(KEYINPUT41), .ZN(new_n616));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  OAI22_X1  g416(.A1(new_n615), .A2(KEYINPUT101), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n549), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(KEYINPUT101), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n616), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n603), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n612), .B(new_n590), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(KEYINPUT10), .ZN(new_n633));
  INV_X1    g432(.A(G230gat), .ZN(new_n634));
  INV_X1    g433(.A(G233gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n632), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n643), .A2(new_n639), .A3(new_n642), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n639), .B2(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND4_X1   g445(.A1(new_n537), .A2(new_n580), .A3(new_n630), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n494), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND3_X1   g449(.A1(new_n647), .A2(new_n497), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n551), .B1(new_n647), .B2(new_n497), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n655), .A3(new_n297), .ZN(new_n656));
  INV_X1    g455(.A(new_n487), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n658), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g458(.A1(new_n647), .A2(new_n488), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT103), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(new_n580), .ZN(new_n664));
  INV_X1    g463(.A(new_n646), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n602), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n537), .A2(new_n629), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G29gat), .A3(new_n466), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n533), .A2(new_n536), .A3(new_n629), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n466), .A2(new_n412), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n451), .A2(new_n455), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n522), .B1(new_n400), .B2(new_n403), .ZN(new_n676));
  INV_X1    g475(.A(new_n523), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT38), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n675), .A2(new_n678), .A3(new_n408), .A4(new_n529), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n417), .B1(new_n506), .B2(new_n508), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n680), .B(new_n513), .C1(new_n506), .C2(new_n503), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n511), .B(new_n681), .C1(new_n449), .C2(new_n450), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n497), .A2(new_n683), .B1(new_n374), .B2(new_n370), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n674), .A2(new_n488), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT105), .B1(new_n685), .B2(new_n487), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n487), .A2(new_n498), .A3(new_n531), .A4(KEYINPUT105), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n480), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT106), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n532), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n479), .B1(new_n692), .B2(new_n687), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n628), .A2(KEYINPUT44), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n692), .A2(new_n687), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n694), .B1(new_n700), .B2(new_n480), .ZN(new_n701));
  AOI211_X1 g500(.A(KEYINPUT106), .B(new_n479), .C1(new_n692), .C2(new_n687), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(KEYINPUT107), .A3(new_n696), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n673), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n666), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n703), .B2(new_n696), .ZN(new_n708));
  INV_X1    g507(.A(new_n696), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n701), .A2(new_n702), .A3(new_n698), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n672), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n666), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(new_n494), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n670), .B1(new_n715), .B2(new_n542), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n667), .A2(G36gat), .A3(new_n412), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n714), .A2(new_n497), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n538), .ZN(G1329gat));
  NOR3_X1   g519(.A1(new_n667), .A2(G43gat), .A3(new_n296), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n705), .A2(new_n487), .A3(new_n706), .ZN(new_n724));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n714), .A2(new_n657), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n727), .B2(G43gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g528(.A1(new_n667), .A2(G50gat), .A3(new_n375), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n705), .A2(new_n375), .A3(new_n706), .ZN(new_n732));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT48), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n707), .A2(new_n713), .A3(new_n488), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n731), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n730), .B1(new_n736), .B2(G50gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(KEYINPUT109), .A3(KEYINPUT48), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n740), .B2(new_n742), .ZN(G1331gat));
  AND4_X1   g542(.A1(new_n664), .A2(new_n703), .A3(new_n630), .A4(new_n665), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n494), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n497), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n657), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n296), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n488), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n580), .A2(new_n602), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n711), .A2(new_n665), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n607), .B1(new_n758), .B2(new_n494), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n629), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n693), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(KEYINPUT51), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n762), .B2(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(new_n761), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n765), .A2(new_n762), .A3(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n466), .A2(new_n646), .A3(G85gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n759), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1336gat));
  AOI21_X1  g571(.A(new_n608), .B1(new_n758), .B2(new_n497), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT51), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n412), .A2(new_n646), .A3(G92gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  INV_X1    g577(.A(new_n776), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n767), .B2(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n777), .A2(new_n778), .B1(new_n773), .B2(new_n780), .ZN(G1337gat));
  XNOR2_X1  g580(.A(KEYINPUT113), .B(G99gat), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n758), .B2(new_n657), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n665), .A2(new_n297), .A3(new_n782), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n768), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n758), .B2(new_n488), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n375), .A2(new_n646), .A3(G106gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n775), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n793));
  INV_X1    g592(.A(new_n790), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n767), .B2(new_n794), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n791), .A2(new_n792), .B1(new_n789), .B2(new_n795), .ZN(G1339gat));
  NOR2_X1   g595(.A1(new_n633), .A2(new_n637), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n638), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n642), .B1(new_n638), .B2(new_n798), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n802), .A2(KEYINPUT55), .B1(new_n639), .B2(new_n642), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n802), .A2(KEYINPUT55), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n580), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n563), .A2(new_n564), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n568), .A2(new_n569), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n576), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n578), .A2(new_n665), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n629), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  AND4_X1   g613(.A1(new_n578), .A2(new_n808), .A3(new_n629), .A4(new_n812), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n603), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n630), .A2(new_n646), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n580), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n376), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n494), .A3(new_n412), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n205), .A3(new_n664), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n475), .A2(new_n477), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n821), .A2(new_n466), .A3(new_n497), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n580), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n824), .A2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n823), .B2(new_n646), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT117), .Z(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(new_n203), .A3(new_n665), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  NOR3_X1   g631(.A1(new_n823), .A2(new_n208), .A3(new_n603), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT118), .Z(new_n834));
  AOI21_X1  g633(.A(G127gat), .B1(new_n826), .B2(new_n602), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n466), .ZN(new_n837));
  INV_X1    g636(.A(new_n825), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n497), .A2(new_n628), .ZN(new_n839));
  XNOR2_X1  g638(.A(KEYINPUT69), .B(G134gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT56), .Z(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n823), .B2(new_n628), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n375), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n807), .A2(new_n803), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n813), .B1(new_n664), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n815), .B1(new_n628), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n602), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n818), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n488), .A2(KEYINPUT57), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n845), .A2(KEYINPUT57), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n657), .A2(new_n466), .A3(new_n497), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n664), .A2(new_n300), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(KEYINPUT58), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n488), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n657), .A3(new_n497), .ZN(new_n860));
  AOI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n580), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n862), .B(new_n863), .Z(G1344gat));
  NAND2_X1  g663(.A1(new_n309), .A2(new_n311), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n860), .A2(new_n866), .A3(new_n665), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n866), .C1(new_n854), .C2(new_n665), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n850), .A2(new_n375), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .B1(new_n821), .B2(new_n851), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n665), .A3(new_n853), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n867), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(G1345gat));
  AOI21_X1  g675(.A(new_n321), .B1(new_n854), .B2(new_n602), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n860), .A2(new_n321), .A3(new_n602), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT121), .Z(G1346gat));
  NAND2_X1  g679(.A1(new_n854), .A2(new_n629), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n322), .B1(new_n881), .B2(KEYINPUT122), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(KEYINPUT122), .B2(new_n881), .ZN(new_n883));
  INV_X1    g682(.A(new_n859), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n322), .A3(new_n487), .A4(new_n839), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n494), .A2(new_n412), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n822), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n220), .A3(new_n664), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n838), .A2(new_n497), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT123), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(KEYINPUT123), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n821), .A2(new_n494), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n580), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n889), .A2(new_n895), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n888), .B2(new_n646), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n221), .A3(new_n665), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1349gat));
  NOR2_X1   g698(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n888), .B2(new_n603), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n240), .A3(new_n602), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n903), .B(new_n904), .Z(G1350gat));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n231), .A3(new_n629), .ZN(new_n906));
  OAI21_X1  g705(.A(G190gat), .B1(new_n888), .B2(new_n628), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n907), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n487), .A2(new_n887), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n821), .A2(new_n375), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n580), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n871), .A2(new_n487), .A3(new_n887), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n580), .A2(G197gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G1352gat));
  AND4_X1   g717(.A1(new_n487), .A2(new_n871), .A3(new_n665), .A4(new_n887), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT126), .B(G204gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n665), .A3(new_n920), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(KEYINPUT62), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(KEYINPUT62), .B2(new_n922), .ZN(G1353gat));
  NAND3_X1  g723(.A1(new_n914), .A2(new_n341), .A3(new_n602), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n916), .A2(new_n602), .ZN(new_n926));
  AND4_X1   g725(.A1(KEYINPUT127), .A2(new_n926), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n927));
  OAI21_X1  g726(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n926), .A2(new_n929), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n927), .B2(new_n930), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n342), .A3(new_n629), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n916), .A2(new_n629), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n342), .ZN(G1355gat));
endmodule


