

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n342), .B(KEYINPUT45), .ZN(n343) );
  XNOR2_X1 U323 ( .A(n344), .B(n343), .ZN(n361) );
  XOR2_X1 U324 ( .A(G29GAT), .B(G134GAT), .Z(n311) );
  XNOR2_X1 U325 ( .A(n295), .B(n294), .ZN(n296) );
  NOR2_X1 U326 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U328 ( .A(KEYINPUT36), .B(n551), .Z(n578) );
  XNOR2_X1 U329 ( .A(n305), .B(n304), .ZN(n551) );
  XNOR2_X1 U330 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U331 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT9), .B(n311), .Z(n291) );
  XOR2_X1 U333 ( .A(G43GAT), .B(G99GAT), .Z(n430) );
  XNOR2_X1 U334 ( .A(n430), .B(G218GAT), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n297) );
  XOR2_X1 U336 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n293) );
  XNOR2_X1 U337 ( .A(G106GAT), .B(G92GAT), .ZN(n292) );
  XOR2_X1 U338 ( .A(n293), .B(n292), .Z(n295) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U340 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n299) );
  XNOR2_X1 U341 ( .A(G162GAT), .B(G85GAT), .ZN(n298) );
  XOR2_X1 U342 ( .A(n299), .B(n298), .Z(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n305) );
  XNOR2_X1 U344 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n302), .B(KEYINPUT7), .ZN(n379) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n303), .B(KEYINPUT75), .ZN(n393) );
  XNOR2_X1 U348 ( .A(n379), .B(n393), .ZN(n304) );
  INV_X1 U349 ( .A(n551), .ZN(n467) );
  XOR2_X1 U350 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n307) );
  XNOR2_X1 U351 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n319) );
  XOR2_X1 U353 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n309) );
  XNOR2_X1 U354 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n315) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G85GAT), .ZN(n310) );
  XOR2_X1 U357 ( .A(n310), .B(G57GAT), .Z(n347) );
  XNOR2_X1 U358 ( .A(n347), .B(n311), .ZN(n313) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U361 ( .A(n315), .B(n314), .Z(n317) );
  XOR2_X1 U362 ( .A(G113GAT), .B(G1GAT), .Z(n378) );
  XOR2_X1 U363 ( .A(KEYINPUT0), .B(G127GAT), .Z(n429) );
  XNOR2_X1 U364 ( .A(n378), .B(n429), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U367 ( .A(G148GAT), .B(G155GAT), .Z(n321) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n323) );
  XNOR2_X1 U371 ( .A(G162GAT), .B(KEYINPUT88), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n417) );
  XNOR2_X1 U374 ( .A(n326), .B(n417), .ZN(n463) );
  XNOR2_X1 U375 ( .A(KEYINPUT94), .B(n463), .ZN(n512) );
  INV_X1 U376 ( .A(KEYINPUT54), .ZN(n411) );
  XNOR2_X1 U377 ( .A(G8GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(KEYINPUT77), .ZN(n396) );
  XOR2_X1 U379 ( .A(KEYINPUT78), .B(G64GAT), .Z(n329) );
  XNOR2_X1 U380 ( .A(G1GAT), .B(G57GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n396), .B(n330), .Z(n332) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G15GAT), .Z(n377) );
  XOR2_X1 U384 ( .A(G71GAT), .B(KEYINPUT13), .Z(n351) );
  XNOR2_X1 U385 ( .A(n377), .B(n351), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U387 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n334) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U391 ( .A(G78GAT), .B(G211GAT), .Z(n338) );
  XNOR2_X1 U392 ( .A(G127GAT), .B(G155GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(KEYINPUT12), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n575) );
  NOR2_X1 U396 ( .A1(n578), .A2(n575), .ZN(n344) );
  INV_X1 U397 ( .A(KEYINPUT114), .ZN(n342) );
  XOR2_X1 U398 ( .A(G64GAT), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n400), .B(n347), .ZN(n360) );
  XOR2_X1 U402 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n349) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G148GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n354), .B(KEYINPUT33), .ZN(n358) );
  XOR2_X1 U409 ( .A(G78GAT), .B(KEYINPUT71), .Z(n356) );
  XNOR2_X1 U410 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n413) );
  XOR2_X1 U412 ( .A(n413), .B(KEYINPUT70), .Z(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n570) );
  NOR2_X1 U415 ( .A1(n361), .A2(n570), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n362), .B(KEYINPUT115), .ZN(n384) );
  XOR2_X1 U417 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n364) );
  XNOR2_X1 U418 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n383) );
  XOR2_X1 U420 ( .A(G141GAT), .B(G36GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G29GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U423 ( .A(KEYINPUT67), .B(G8GAT), .Z(n368) );
  XNOR2_X1 U424 ( .A(G169GAT), .B(G197GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U426 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U427 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n372) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT29), .B(n373), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n381) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U435 ( .A(n383), .B(n382), .Z(n566) );
  INV_X1 U436 ( .A(n566), .ZN(n542) );
  NOR2_X1 U437 ( .A1(n384), .A2(n542), .ZN(n391) );
  XNOR2_X1 U438 ( .A(KEYINPUT41), .B(n570), .ZN(n559) );
  NOR2_X1 U439 ( .A1(n559), .A2(n566), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  XNOR2_X1 U441 ( .A(KEYINPUT113), .B(n386), .ZN(n388) );
  INV_X1 U442 ( .A(n575), .ZN(n549) );
  NOR2_X1 U443 ( .A1(n551), .A2(n549), .ZN(n387) );
  AND2_X1 U444 ( .A1(n388), .A2(n387), .ZN(n389) );
  XOR2_X1 U445 ( .A(n389), .B(KEYINPUT47), .Z(n390) );
  XNOR2_X1 U446 ( .A(n392), .B(KEYINPUT48), .ZN(n525) );
  XOR2_X1 U447 ( .A(KEYINPUT95), .B(n393), .Z(n395) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n402) );
  XOR2_X1 U451 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n399) );
  XNOR2_X1 U452 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n434) );
  XNOR2_X1 U454 ( .A(n434), .B(n400), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n408) );
  XNOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT85), .ZN(n404) );
  XOR2_X1 U458 ( .A(n404), .B(KEYINPUT21), .Z(n406) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n414) );
  INV_X1 U461 ( .A(n414), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n516) );
  XNOR2_X1 U463 ( .A(n516), .B(KEYINPUT121), .ZN(n409) );
  NOR2_X1 U464 ( .A1(n525), .A2(n409), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X2 U466 ( .A1(n512), .A2(n412), .ZN(n565) );
  XOR2_X1 U467 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n416) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n426) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XOR2_X1 U472 ( .A(G204GAT), .B(KEYINPUT89), .Z(n420) );
  XNOR2_X1 U473 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U475 ( .A(G50GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n457) );
  NAND2_X1 U479 ( .A1(n565), .A2(n457), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n427), .B(KEYINPUT55), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n428), .B(KEYINPUT122), .ZN(n448) );
  XOR2_X1 U482 ( .A(G190GAT), .B(G134GAT), .Z(n432) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U485 ( .A(n433), .B(G71GAT), .Z(n439) );
  XOR2_X1 U486 ( .A(n434), .B(G15GAT), .Z(n436) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(G113GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n447) );
  XOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n441) );
  XNOR2_X1 U492 ( .A(G176GAT), .B(G183GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U494 ( .A(G120GAT), .B(KEYINPUT20), .Z(n443) );
  XNOR2_X1 U495 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U497 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n528) );
  NAND2_X1 U499 ( .A1(n448), .A2(n528), .ZN(n562) );
  NOR2_X1 U500 ( .A1(n467), .A2(n562), .ZN(n451) );
  XNOR2_X1 U501 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n516), .B(KEYINPUT27), .ZN(n460) );
  NAND2_X1 U503 ( .A1(n512), .A2(n460), .ZN(n524) );
  NOR2_X1 U504 ( .A1(n528), .A2(n524), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n457), .B(KEYINPUT28), .ZN(n527) );
  NAND2_X1 U506 ( .A1(n452), .A2(n527), .ZN(n453) );
  XOR2_X1 U507 ( .A(KEYINPUT96), .B(n453), .Z(n466) );
  NAND2_X1 U508 ( .A1(n528), .A2(n516), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n454), .A2(n457), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(KEYINPUT98), .ZN(n462) );
  NOR2_X1 U512 ( .A1(n457), .A2(n528), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT97), .B(n458), .Z(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT26), .B(n459), .Z(n541) );
  INV_X1 U515 ( .A(n541), .ZN(n564) );
  AND2_X1 U516 ( .A1(n564), .A2(n460), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n484) );
  XOR2_X1 U520 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n469) );
  NAND2_X1 U521 ( .A1(n549), .A2(n467), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n484), .A2(n470), .ZN(n498) );
  NOR2_X1 U524 ( .A1(n566), .A2(n570), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT73), .B(n471), .Z(n487) );
  NAND2_X1 U526 ( .A1(n498), .A2(n487), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT99), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n482), .A2(n512), .ZN(n476) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n474) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n482), .A2(n516), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT102), .ZN(n478) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n478), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U537 ( .A1(n482), .A2(n528), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  INV_X1 U540 ( .A(n527), .ZN(n520) );
  NAND2_X1 U541 ( .A1(n482), .A2(n520), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NOR2_X1 U544 ( .A1(n578), .A2(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n575), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n486), .ZN(n511) );
  NAND2_X1 U547 ( .A1(n511), .A2(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n488), .Z(n495) );
  NAND2_X1 U549 ( .A1(n512), .A2(n495), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n516), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n528), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  XOR2_X1 U557 ( .A(G50GAT), .B(KEYINPUT105), .Z(n497) );
  NAND2_X1 U558 ( .A1(n520), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  NOR2_X1 U560 ( .A1(n559), .A2(n542), .ZN(n510) );
  AND2_X1 U561 ( .A1(n498), .A2(n510), .ZN(n505) );
  NAND2_X1 U562 ( .A1(n505), .A2(n512), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n500) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n505), .A2(n516), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n528), .A2(n505), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U572 ( .A1(n505), .A2(n520), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT108), .Z(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n514) );
  AND2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n512), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n528), .A2(n521), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT112), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT116), .B(n526), .Z(n540) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n540), .A2(n529), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n542), .A2(n536), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n532) );
  INV_X1 U596 ( .A(n559), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n536), .A2(n544), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NAND2_X1 U600 ( .A1(n549), .A2(n536), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U604 ( .A1(n536), .A2(n551), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U611 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n562), .A2(n566), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT123), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n559), .A2(n562), .ZN(n560) );
  XOR2_X1 U627 ( .A(n561), .B(n560), .Z(G1349GAT) );
  NOR2_X1 U628 ( .A1(n575), .A2(n562), .ZN(n563) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n577), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

