//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n204), .A2(new_n205), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n216), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n202), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n211), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n225), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n220), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n209), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n254), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n208), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n262), .B(new_n267), .C1(G50), .C2(new_n263), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n273), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n291), .A3(G274), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(G226), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n272), .B1(new_n299), .B2(G190), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n272), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n298), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n300), .B(new_n305), .C1(new_n301), .C2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n268), .C1(G179), .C2(new_n298), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n281), .B2(G20), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n277), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT74), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n202), .A2(new_n203), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n217), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n259), .A2(G159), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n203), .B1(new_n315), .B2(new_n316), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n328), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n333), .A3(new_n254), .ZN(new_n334));
  INV_X1    g0134(.A(new_n265), .ZN(new_n335));
  INV_X1    g0135(.A(new_n256), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n266), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n335), .A2(new_n337), .B1(new_n263), .B2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT75), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n292), .B1(new_n227), .B2(new_n295), .ZN(new_n341));
  INV_X1    g0141(.A(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n283), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G226), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n345), .C1(new_n318), .C2(new_n319), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n291), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n347), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n273), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n296), .A2(G232), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n292), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n310), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n349), .A2(new_n340), .A3(new_n350), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n334), .A2(new_n339), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT18), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT76), .B1(new_n355), .B2(G190), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT76), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(new_n364), .A3(new_n306), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n334), .A3(new_n339), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n209), .A2(G33), .A3(G77), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n203), .A2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n218), .B2(new_n260), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n254), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT11), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT11), .B(new_n254), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(KEYINPUT71), .A3(new_n379), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n208), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n386), .B(KEYINPUT12), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n384), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n344), .A2(new_n342), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n227), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n318), .C2(new_n319), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n273), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n291), .A2(G238), .A3(new_n294), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n292), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n291), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n292), .A2(new_n399), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT13), .ZN(new_n404));
  OAI21_X1  g0204(.A(G200), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(new_n400), .A3(new_n392), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT13), .B1(new_n402), .B2(new_n403), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(G190), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n391), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n401), .B2(new_n404), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT73), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n310), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n406), .A2(G179), .A3(new_n407), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n410), .B1(new_n421), .B2(new_n391), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n256), .B(KEYINPUT68), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n260), .ZN(new_n425));
  INV_X1    g0225(.A(G87), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT15), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT15), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n431), .A2(new_n257), .B1(new_n209), .B2(new_n284), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n254), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n284), .B1(new_n208), .B2(G20), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n265), .A2(new_n434), .B1(new_n284), .B2(new_n264), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n278), .A2(G232), .B1(new_n320), .B2(G107), .ZN(new_n437));
  INV_X1    g0237(.A(G238), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n282), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n273), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n293), .B1(G244), .B2(new_n296), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n350), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n310), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n436), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(new_n435), .C1(new_n306), .C2(new_n443), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n362), .B1(new_n440), .B2(new_n441), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n422), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n313), .A2(new_n369), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n208), .A2(G45), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n273), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n455), .ZN(new_n458));
  INV_X1    g0258(.A(G274), .ZN(new_n459));
  INV_X1    g0259(.A(new_n220), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n290), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n457), .A2(G270), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(G257), .B(new_n342), .C1(new_n318), .C2(new_n319), .ZN(new_n463));
  INV_X1    g0263(.A(G303), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n281), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n281), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G190), .B(new_n462), .C1(new_n470), .C2(new_n291), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n264), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n254), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n263), .C1(G1), .C2(new_n275), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(new_n472), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n253), .A2(new_n220), .B1(G20), .B2(new_n472), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(G33), .B2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n275), .A2(G97), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT20), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT20), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n476), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n471), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n468), .A2(new_n469), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n320), .A2(G303), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n490), .A2(new_n463), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n273), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n362), .B1(new_n493), .B2(new_n462), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n453), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n462), .B1(new_n470), .B2(new_n291), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n487), .A4(new_n471), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n291), .B1(new_n489), .B2(new_n491), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n457), .A2(G270), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n458), .A2(new_n461), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(G169), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n500), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n485), .A2(new_n486), .ZN(new_n507));
  INV_X1    g0307(.A(new_n476), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n496), .A3(KEYINPUT21), .A4(G169), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n496), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n509), .A3(new_n513), .A4(G179), .ZN(new_n514));
  OAI211_X1 g0314(.A(G179), .B(new_n462), .C1(new_n470), .C2(new_n291), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT82), .B1(new_n515), .B2(new_n487), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n499), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n263), .A2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(new_n475), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(G97), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n259), .A2(G77), .ZN(new_n523));
  INV_X1    g0323(.A(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n523), .B1(new_n529), .B2(new_n209), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n524), .B1(new_n315), .B2(new_n316), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n254), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT77), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT7), .B1(new_n320), .B2(new_n209), .ZN(new_n534));
  INV_X1    g0334(.A(new_n316), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n474), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n522), .B1(new_n533), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G283), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n547));
  OAI211_X1 g0347(.A(G244), .B(new_n342), .C1(new_n318), .C2(new_n319), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT4), .B1(new_n278), .B2(G244), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n273), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n457), .A2(G257), .B1(new_n458), .B2(new_n461), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n350), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G169), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT78), .B1(new_n545), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n542), .A2(new_n543), .ZN(new_n558));
  AOI211_X1 g0358(.A(KEYINPUT77), .B(new_n474), .C1(new_n536), .C2(new_n541), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n521), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g0361(.A(G169), .B1(new_n552), .B2(new_n553), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n350), .B2(new_n555), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n552), .A2(new_n553), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n555), .A2(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n545), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n291), .A2(G250), .A3(new_n454), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n291), .A2(G274), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n454), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n281), .A2(G244), .A3(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(G238), .B(new_n342), .C1(new_n318), .C2(new_n319), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n576), .B2(new_n273), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G190), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n362), .B2(new_n577), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n520), .A2(G87), .ZN(new_n581));
  NAND3_X1  g0381(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n209), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n538), .A2(new_n426), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n209), .B(G68), .C1(new_n318), .C2(new_n319), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n257), .B2(new_n228), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n254), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n430), .A2(new_n263), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT79), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT79), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n594), .B(new_n591), .C1(new_n589), .C2(new_n254), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n581), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n580), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n577), .A2(G169), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n350), .B2(new_n577), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n520), .A2(new_n430), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n593), .B2(new_n595), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n604));
  OAI211_X1 g0404(.A(G250), .B(new_n342), .C1(new_n318), .C2(new_n319), .ZN(new_n605));
  INV_X1    g0405(.A(G294), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n604), .B(new_n605), .C1(new_n275), .C2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n273), .B1(new_n457), .B2(G264), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n503), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n310), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n350), .A3(new_n503), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT23), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n524), .A3(G20), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n612), .A2(new_n614), .A3(new_n615), .A4(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n209), .B(G87), .C1(new_n318), .C2(new_n319), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT22), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n281), .A2(new_n623), .A3(new_n209), .A4(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT24), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT24), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n620), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n474), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n475), .A2(new_n524), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n263), .A2(G107), .ZN(new_n632));
  XNOR2_X1  g0432(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n610), .B(new_n611), .C1(new_n630), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n629), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n628), .B1(new_n620), .B2(new_n625), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n254), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n608), .A2(G190), .A3(new_n503), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n609), .A2(G200), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n640), .A2(new_n635), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n598), .A2(new_n603), .A3(new_n637), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n518), .A2(new_n569), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n452), .A2(new_n645), .ZN(G372));
  INV_X1    g0446(.A(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n359), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n421), .A2(new_n391), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n410), .B2(new_n445), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(new_n368), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n308), .A2(new_n309), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n312), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n511), .A2(new_n517), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n637), .A2(KEYINPUT88), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n637), .A2(KEYINPUT88), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n590), .A2(new_n592), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n594), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n590), .A2(KEYINPUT79), .A3(new_n592), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT86), .B1(new_n663), .B2(new_n581), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n581), .B(KEYINPUT86), .C1(new_n593), .C2(new_n595), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n580), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n603), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT86), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n596), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n579), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n577), .A2(new_n350), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(G169), .B2(new_n577), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n663), .B2(new_n601), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT87), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n643), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n569), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n659), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT89), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n545), .A2(new_n556), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI211_X1 g0484(.A(KEYINPUT26), .B(new_n684), .C1(new_n669), .C2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n598), .A2(new_n603), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n557), .B2(new_n564), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n603), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n682), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n677), .A2(new_n688), .A3(new_n683), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n597), .A2(new_n580), .B1(new_n600), .B2(new_n602), .ZN(new_n692));
  INV_X1    g0492(.A(new_n564), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n675), .B1(new_n695), .B2(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n696), .A3(KEYINPUT89), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n681), .B1(new_n690), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n452), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n654), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT90), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n509), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n499), .A2(new_n511), .A3(new_n517), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n655), .B2(new_n708), .ZN(new_n710));
  INV_X1    g0510(.A(new_n637), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n707), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n640), .A2(new_n635), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n707), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n637), .A3(new_n643), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(G330), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n511), .A2(new_n517), .ZN(new_n718));
  INV_X1    g0518(.A(new_n707), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n637), .A3(new_n643), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n658), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n656), .A3(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n717), .A2(new_n724), .ZN(G399));
  NOR2_X1   g0525(.A1(new_n213), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n584), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n219), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n727), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n691), .A2(new_n696), .A3(KEYINPUT89), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT89), .B1(new_n691), .B2(new_n696), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n680), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n719), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n688), .B1(new_n677), .B2(new_n683), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n603), .B1(new_n695), .B2(KEYINPUT26), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n679), .B(new_n677), .C1(new_n718), .C2(new_n711), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n719), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n577), .A2(new_n608), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n515), .A2(new_n746), .A3(new_n565), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n577), .A2(G179), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n496), .A3(new_n565), .A4(new_n609), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n555), .A2(new_n577), .A3(new_n608), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n752), .B2(new_n515), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n707), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n499), .A2(new_n511), .A3(new_n517), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n557), .A2(new_n564), .A3(new_n568), .ZN(new_n758));
  INV_X1    g0558(.A(new_n644), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n719), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n756), .B1(new_n760), .B2(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n751), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n747), .A2(new_n748), .ZN(new_n763));
  OAI211_X1 g0563(.A(KEYINPUT31), .B(new_n707), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(G330), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n745), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n732), .B1(new_n767), .B2(G1), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT91), .ZN(G364));
  AND2_X1   g0569(.A1(new_n209), .A2(G13), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n208), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n726), .A2(KEYINPUT92), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT92), .B1(new_n726), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n220), .B1(G20), .B2(new_n310), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n209), .A2(new_n306), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n350), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n209), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n779), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n320), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n782), .B(new_n786), .C1(G329), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n362), .A2(G179), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n778), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G303), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n783), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G283), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n209), .B1(new_n787), .B2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n306), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(G294), .B1(G326), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n802), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  OAI211_X1 g0607(.A(new_n799), .B(new_n804), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n780), .ZN(new_n809));
  INV_X1    g0609(.A(new_n784), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G58), .A2(new_n809), .B1(new_n810), .B2(G77), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(KEYINPUT93), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G87), .B2(new_n794), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(G107), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n789), .A2(G159), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT32), .ZN(new_n816));
  INV_X1    g0616(.A(new_n803), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n806), .A2(new_n203), .B1(new_n817), .B2(new_n218), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n800), .A2(new_n228), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n320), .B(new_n820), .C1(new_n811), .C2(KEYINPUT93), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n813), .A2(new_n814), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n777), .B1(new_n808), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n776), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n219), .A2(new_n288), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n213), .A2(new_n281), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n248), .C2(new_n288), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n213), .A2(new_n320), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G355), .B1(new_n472), .B2(new_n213), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n775), .B(new_n823), .C1(new_n827), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n826), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n710), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n710), .A2(G330), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n775), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n710), .A2(G330), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n775), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n436), .A2(new_n707), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n447), .B2(new_n448), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n445), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n445), .A2(new_n707), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n698), .B2(new_n707), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n450), .A2(new_n719), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n698), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n841), .B1(new_n850), .B2(new_n766), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n766), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n776), .A2(new_n824), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(G77), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n798), .A2(G68), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n218), .B2(new_n793), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT95), .Z(new_n858));
  AOI21_X1  g0658(.A(new_n320), .B1(new_n789), .B2(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n202), .B2(new_n800), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n809), .B1(new_n810), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n861), .B1(new_n806), .B2(new_n258), .C1(new_n862), .C2(new_n817), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT34), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n820), .B1(new_n803), .B2(G303), .ZN(new_n867));
  INV_X1    g0667(.A(G283), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n806), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n780), .A2(new_n606), .B1(new_n784), .B2(new_n472), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n281), .B(new_n870), .C1(G311), .C2(new_n789), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n798), .A2(G87), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n871), .B(new_n872), .C1(new_n524), .C2(new_n793), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n858), .A2(new_n866), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n855), .B1(new_n874), .B2(new_n776), .ZN(new_n875));
  INV_X1    g0675(.A(new_n847), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n825), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n852), .A2(new_n877), .ZN(G384));
  OR2_X1    g0678(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(G116), .A3(new_n221), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  OAI211_X1 g0682(.A(new_n219), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n203), .A2(G50), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT96), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n208), .B(G13), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n745), .A2(new_n699), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n653), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n328), .B1(new_n323), .B2(G68), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n474), .B1(new_n890), .B2(KEYINPUT16), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n324), .A2(new_n329), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n331), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n339), .ZN(new_n895));
  INV_X1    g0695(.A(new_n705), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n360), .B2(new_n368), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n357), .A2(new_n358), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n897), .A3(new_n367), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n366), .A2(new_n334), .A3(new_n339), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n359), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n705), .B1(new_n334), .B2(new_n339), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n901), .A2(KEYINPUT37), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n898), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n897), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT17), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n367), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n648), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n338), .B1(new_n891), .B2(new_n893), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n367), .B1(new_n913), .B2(new_n705), .ZN(new_n914));
  INV_X1    g0714(.A(new_n899), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n903), .A2(new_n905), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n908), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT98), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n338), .B1(new_n891), .B2(new_n333), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n705), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n367), .B1(new_n915), .B2(new_n924), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT37), .B(new_n925), .C1(new_n926), .C2(new_n904), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT37), .B1(new_n904), .B2(KEYINPUT98), .ZN(new_n928));
  INV_X1    g0728(.A(new_n904), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n903), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT99), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n904), .B1(new_n648), .B2(new_n911), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT99), .B1(new_n927), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n907), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n922), .B1(new_n937), .B2(new_n921), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n649), .A2(new_n707), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n846), .B1(new_n698), .B2(new_n849), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n907), .B1(new_n898), .B2(new_n906), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n936), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n421), .A2(new_n391), .A3(new_n707), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT97), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n391), .A2(new_n707), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n422), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n383), .A2(new_n390), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n948), .A2(new_n382), .A3(new_n408), .A4(new_n405), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n419), .B1(new_n416), .B2(new_n412), .ZN(new_n950));
  INV_X1    g0750(.A(new_n391), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n949), .B(new_n946), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(KEYINPUT97), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n944), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n941), .A2(new_n943), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n648), .A2(new_n705), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n940), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n889), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n952), .A2(KEYINPUT97), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n649), .A2(new_n945), .A3(new_n949), .A4(new_n946), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n847), .B1(new_n962), .B2(new_n944), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n754), .A2(KEYINPUT100), .A3(KEYINPUT31), .A4(new_n707), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT100), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n764), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n963), .B(KEYINPUT40), .C1(new_n761), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n964), .A2(new_n966), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT31), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n645), .B2(new_n719), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n972), .B2(new_n756), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n943), .A3(new_n963), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT40), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n969), .A2(new_n937), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n760), .A2(KEYINPUT31), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n967), .B1(new_n978), .B2(new_n755), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n977), .B1(new_n699), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n452), .A3(new_n973), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(G330), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n959), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n208), .B2(new_n770), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n959), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n887), .B1(new_n984), .B2(new_n985), .ZN(G367));
  INV_X1    g0786(.A(new_n829), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n827), .B1(new_n212), .B2(new_n431), .C1(new_n987), .C2(new_n243), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n841), .A2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n780), .A2(new_n258), .B1(new_n784), .B2(new_n218), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n320), .B(new_n990), .C1(G137), .C2(new_n789), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n798), .A2(G77), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n202), .C2(new_n793), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n800), .A2(new_n203), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n803), .B2(G143), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n806), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n793), .A2(new_n472), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n798), .A2(G97), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n806), .A2(new_n606), .B1(new_n817), .B2(new_n785), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G107), .B2(new_n801), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n281), .B1(new_n809), .B2(G303), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n810), .B1(new_n789), .B2(G317), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n993), .A2(new_n997), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  NAND3_X1  g0807(.A1(new_n671), .A2(new_n665), .A3(new_n707), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n603), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n677), .B2(new_n1008), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n989), .B1(new_n777), .B2(new_n1007), .C1(new_n1011), .C2(new_n835), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT105), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n718), .A2(new_n719), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1014), .A2(new_n715), .A3(new_n712), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT103), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(KEYINPUT103), .A3(new_n715), .A4(new_n712), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n720), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT104), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n837), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT104), .B1(new_n710), .B2(G330), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1022), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1024), .A2(new_n720), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n745), .A2(new_n1013), .A3(new_n766), .A4(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1026), .A2(new_n737), .A3(new_n744), .A4(new_n766), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT105), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n758), .B1(new_n545), .B2(new_n719), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n683), .A2(new_n707), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n724), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT44), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n724), .B2(new_n1032), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n723), .A2(KEYINPUT44), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1035), .A2(new_n717), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n717), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1027), .A2(new_n1029), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n767), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n726), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n772), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1030), .A2(KEYINPUT101), .A3(new_n1031), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT101), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n711), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n693), .A2(new_n694), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n707), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n720), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1032), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT42), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT102), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT102), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1048), .B(new_n1060), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1062), .A2(new_n1063), .B1(new_n717), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1059), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1065), .A2(new_n717), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1012), .B1(new_n1047), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT106), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(KEYINPUT106), .B(new_n1012), .C1(new_n1047), .C2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G387));
  NAND2_X1  g0879(.A1(new_n1026), .A2(new_n772), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n780), .A2(new_n218), .B1(new_n788), .B2(new_n258), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n320), .B(new_n1081), .C1(G68), .C2(new_n810), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n996), .A2(new_n817), .B1(new_n806), .B2(new_n256), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n431), .A2(new_n800), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n794), .A2(G77), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1000), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n281), .B1(new_n789), .B2(G326), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n793), .A2(new_n606), .B1(new_n868), .B2(new_n800), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n809), .B1(new_n810), .B2(G303), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n806), .B2(new_n785), .C1(new_n781), .C2(new_n817), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1088), .B1(new_n472), .B2(new_n797), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n776), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n712), .A2(new_n715), .A3(new_n826), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n728), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n831), .A2(new_n1101), .B1(new_n524), .B2(new_n213), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n423), .A2(new_n218), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT50), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n288), .B1(new_n203), .B2(new_n284), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1104), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n829), .B1(new_n240), .B2(new_n288), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1102), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(KEYINPUT107), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT107), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n827), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1099), .A2(new_n841), .A3(new_n1100), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n726), .B1(new_n767), .B2(new_n1026), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1080), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(G393));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1042), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1043), .A2(new_n726), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1042), .A2(new_n772), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT108), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1065), .A2(new_n826), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n320), .B1(new_n784), .B2(new_n606), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n806), .A2(new_n464), .B1(new_n800), .B2(new_n472), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G322), .C2(new_n789), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n814), .C1(new_n868), .C2(new_n793), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n809), .A2(G311), .B1(G317), .B2(new_n803), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n872), .B1(new_n203), .B2(new_n793), .C1(new_n424), .C2(new_n784), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n806), .A2(new_n218), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n320), .B(new_n1128), .C1(G143), .C2(new_n789), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n817), .A2(new_n258), .B1(new_n780), .B2(new_n996), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT51), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n800), .A2(new_n284), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1124), .A2(new_n1126), .B1(new_n1127), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n776), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n829), .A2(new_n251), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1139), .B(new_n827), .C1(new_n228), .C2(new_n212), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1120), .A2(new_n841), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1118), .A2(new_n1119), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1119), .B1(new_n1118), .B2(new_n1141), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1116), .A2(new_n1117), .B1(new_n1142), .B2(new_n1143), .ZN(G390));
  OAI211_X1 g0944(.A(G330), .B(new_n876), .C1(new_n761), .C2(new_n765), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n954), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n939), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n937), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n844), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n846), .B1(new_n743), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1152), .B2(new_n954), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n938), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n939), .B1(new_n941), .B2(new_n954), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT109), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(KEYINPUT109), .B(new_n939), .C1(new_n941), .C2(new_n954), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1148), .B(new_n1154), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n849), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n845), .B1(new_n735), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1149), .B1(new_n1162), .B2(new_n1146), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n938), .B1(new_n1163), .B2(KEYINPUT109), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1153), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n954), .A2(new_n876), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n979), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(G330), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1160), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n973), .A2(G330), .A3(new_n452), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT110), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT110), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n973), .A2(new_n1173), .A3(new_n452), .A4(G330), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n654), .B(new_n1175), .C1(new_n745), .C2(new_n699), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1152), .A2(new_n1147), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n973), .A2(G330), .A3(new_n876), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1146), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1169), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1177), .A2(new_n1179), .B1(new_n1181), .B2(new_n941), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1160), .B(new_n1183), .C1(new_n1166), .C2(new_n1169), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n726), .A3(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1160), .B(new_n772), .C1(new_n1166), .C2(new_n1169), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT112), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n841), .B1(new_n336), .B2(new_n854), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n798), .A2(G50), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT54), .B(G143), .Z(new_n1192));
  AOI21_X1  g0992(.A(new_n320), .B1(new_n810), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G132), .A2(new_n809), .B1(new_n789), .B2(G125), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n805), .A2(G137), .B1(new_n803), .B2(G128), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n996), .C2(new_n800), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n793), .A2(new_n258), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1135), .B1(new_n806), .B2(new_n524), .C1(new_n868), .C2(new_n817), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n780), .A2(new_n472), .B1(new_n788), .B2(new_n606), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n281), .B(new_n1202), .C1(G97), .C2(new_n810), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n856), .C1(new_n426), .C2(new_n793), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1197), .A2(new_n1200), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1190), .B1(new_n1205), .B2(new_n776), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n938), .B2(new_n825), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1188), .A2(new_n1189), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1189), .B1(new_n1188), .B2(new_n1207), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1187), .B1(new_n1208), .B2(new_n1209), .ZN(G378));
  NAND2_X1  g1010(.A1(new_n268), .A2(new_n896), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n313), .A2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n308), .A2(new_n309), .A3(new_n312), .A4(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n976), .B2(G330), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1168), .A2(new_n937), .A3(KEYINPUT40), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n963), .B1(new_n761), .B2(new_n967), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n908), .A2(new_n920), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n975), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AND4_X1   g1025(.A1(G330), .A2(new_n1222), .A3(new_n1225), .A4(new_n1220), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n957), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(G330), .A3(new_n1225), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1220), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n938), .A2(new_n939), .B1(new_n648), .B2(new_n705), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1222), .A2(new_n1225), .A3(new_n1220), .A4(G330), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n955), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n772), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n281), .A2(G41), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G50), .B(new_n1236), .C1(new_n275), .C2(new_n287), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT113), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1236), .B1(new_n524), .B2(new_n780), .C1(new_n868), .C2(new_n788), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n994), .B(new_n1239), .C1(G116), .C2(new_n803), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n810), .A2(new_n430), .B1(G97), .B2(new_n805), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT114), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n798), .A2(G58), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1086), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT58), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1238), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n809), .A2(G128), .B1(G125), .B2(new_n803), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n258), .B2(new_n800), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n810), .A2(G137), .B1(G132), .B2(new_n805), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT115), .Z(new_n1250));
  AOI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n794), .C2(new_n1192), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT116), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  AOI211_X1 g1053(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n996), .C2(new_n797), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1246), .B1(new_n1245), .B2(new_n1244), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n776), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n775), .B1(new_n218), .B2(new_n853), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n1220), .C2(new_n825), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1235), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1176), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1186), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1234), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT117), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1227), .A2(new_n1233), .A3(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n958), .A2(KEYINPUT117), .A3(new_n1232), .A4(new_n1230), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1268), .A2(KEYINPUT57), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n727), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1261), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(G375));
  NOR2_X1   g1073(.A1(new_n954), .A2(new_n825), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1084), .B1(new_n805), .B2(G116), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n606), .B2(new_n817), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n794), .A2(G97), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n281), .B1(new_n809), .B2(G283), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G107), .A2(new_n810), .B1(new_n789), .B2(G303), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n992), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n794), .A2(G159), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n320), .B1(new_n810), .B2(G150), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G137), .A2(new_n809), .B1(new_n789), .B2(G128), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1243), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1192), .A2(new_n805), .B1(G132), .B2(new_n803), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n218), .B2(new_n800), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1276), .A2(new_n1280), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n776), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n841), .C1(G68), .C2(new_n854), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1182), .A2(new_n771), .B1(new_n1274), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1183), .A2(new_n1045), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1292), .A2(KEYINPUT118), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT118), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1291), .B1(new_n1294), .B2(new_n1295), .ZN(G381));
  OR2_X1    g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G381), .A2(new_n1297), .A3(G384), .A4(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1078), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT119), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(G375), .A2(G378), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1298), .A2(KEYINPUT119), .A3(new_n1078), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(G407));
  NAND2_X1  g1104(.A1(new_n706), .A2(G213), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(KEYINPUT120), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G407), .A2(G213), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT121), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(G407), .A2(KEYINPUT121), .A3(G213), .A4(new_n1307), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G409));
  XNOR2_X1  g1112(.A(G393), .B(G396), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G390), .B(new_n1012), .C1(new_n1047), .C2(new_n1073), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G390), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1076), .A2(new_n1077), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1076), .A2(KEYINPUT124), .A3(new_n1077), .A4(new_n1316), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1313), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1074), .A2(new_n1316), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1314), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1319), .A2(new_n1320), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1293), .B1(new_n1183), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1176), .A2(new_n1182), .A3(KEYINPUT60), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n726), .A3(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1329));
  AND2_X1   g1129(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1328), .B(new_n1291), .C1(new_n1329), .C2(new_n1330), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1328), .A2(new_n1291), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1330), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1306), .A2(G2897), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1305), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(G2897), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1268), .A2(new_n772), .A3(new_n1269), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1260), .ZN(new_n1340));
  AOI22_X1  g1140(.A1(new_n1186), .A2(new_n1262), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1341), .B2(new_n1046), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(G378), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1343), .B1(G378), .B2(new_n1272), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1338), .B1(new_n1344), .B2(new_n1306), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1263), .A2(new_n1270), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1346), .B(new_n726), .C1(KEYINPUT57), .C2(new_n1341), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1261), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(G378), .A3(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1263), .A2(new_n1046), .A3(new_n1234), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1340), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1209), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1188), .A2(new_n1189), .A3(new_n1207), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1352), .A2(new_n1355), .A3(new_n1187), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1349), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT62), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1333), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1305), .A4(new_n1359), .ZN(new_n1360));
  XOR2_X1   g1160(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1361));
  NAND3_X1  g1161(.A1(new_n1345), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI211_X1 g1162(.A(new_n1306), .B(new_n1333), .C1(new_n1349), .C2(new_n1356), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1363), .A2(new_n1358), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1324), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT123), .B1(new_n1357), .B2(new_n1305), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT123), .ZN(new_n1367));
  AOI211_X1 g1167(.A(new_n1367), .B(new_n1336), .C1(new_n1349), .C2(new_n1356), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1338), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT63), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1357), .A2(new_n1370), .A3(new_n1305), .A4(new_n1359), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1371), .B1(new_n1363), .B2(new_n1370), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT125), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1373), .B1(new_n1324), .B2(KEYINPUT61), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1315), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1375), .A2(new_n1320), .A3(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1323), .A2(new_n1321), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT61), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1379), .A2(KEYINPUT125), .A3(new_n1380), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1369), .A2(new_n1372), .A3(new_n1374), .A4(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1365), .A2(new_n1382), .ZN(G405));
  NAND3_X1  g1183(.A1(new_n1379), .A2(KEYINPUT127), .A3(new_n1349), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1349), .A2(KEYINPUT127), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1324), .A2(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1384), .A2(new_n1386), .ZN(new_n1387));
  OR2_X1    g1187(.A1(new_n1272), .A2(G378), .ZN(new_n1388));
  XNOR2_X1  g1188(.A(new_n1388), .B(new_n1359), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1387), .A2(new_n1389), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1388), .B(new_n1333), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1391), .A2(new_n1384), .A3(new_n1386), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1390), .A2(new_n1392), .ZN(G402));
endmodule


