//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT91), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n213), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n211), .A2(KEYINPUT91), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(KEYINPUT91), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n211), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n213), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n224), .A2(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(KEYINPUT90), .A3(new_n213), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  AOI21_X1  g035(.A(G1gat), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n222), .B(new_n229), .C1(new_n238), .C2(new_n239), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(KEYINPUT96), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT94), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT96), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n248), .A3(new_n240), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n222), .A2(KEYINPUT17), .A3(new_n229), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n214), .A2(new_n215), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n209), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n255), .B2(new_n228), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n251), .B(new_n256), .C1(new_n238), .C2(new_n239), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n241), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT97), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n245), .A3(new_n241), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n250), .A2(new_n258), .A3(KEYINPUT97), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G141gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G197gat), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT11), .B(G169gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT89), .Z(new_n272));
  INV_X1    g071(.A(new_n259), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n264), .A2(new_n271), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n266), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276));
  INV_X1    g075(.A(G228gat), .ZN(new_n277));
  INV_X1    g076(.A(G233gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G211gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT22), .B1(new_n286), .B2(G218gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G218gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n283), .B2(new_n285), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n288), .B(new_n280), .C1(new_n292), .C2(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n297), .A2(new_n299), .B1(KEYINPUT2), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n303), .A2(new_n307), .A3(new_n310), .A4(new_n304), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n301), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n301), .A2(new_n300), .A3(new_n307), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n295), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n294), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n313), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n290), .B2(new_n293), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n279), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n279), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT81), .B(new_n318), .C1(new_n319), .C2(KEYINPUT3), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n314), .A2(new_n315), .ZN(new_n328));
  INV_X1    g127(.A(new_n293), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT72), .B(G211gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n291), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n280), .B1(new_n332), .B2(new_n288), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n327), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g134(.A(KEYINPUT82), .B(new_n294), .C1(new_n314), .C2(new_n315), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n321), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(G22gat), .B1(new_n338), .B2(KEYINPUT83), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n340), .B(new_n321), .C1(new_n326), .C2(new_n337), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n276), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n321), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n295), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT81), .B1(new_n344), .B2(new_n318), .ZN(new_n345));
  INV_X1    g144(.A(new_n325), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n279), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n316), .B(new_n327), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(KEYINPUT83), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT84), .A4(G22gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n349), .A2(G22gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354));
  INV_X1    g153(.A(G50gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n349), .A2(G22gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n358), .B1(new_n361), .B2(new_n353), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372));
  INV_X1    g171(.A(G113gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G120gat), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(G113gat), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n371), .B(new_n372), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378));
  INV_X1    g177(.A(G127gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G134gat), .ZN(new_n380));
  INV_X1    g179(.A(G134gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(G127gat), .ZN(new_n382));
  OAI22_X1  g181(.A1(new_n378), .A2(KEYINPUT1), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT77), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n318), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n314), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n377), .A2(new_n383), .A3(KEYINPUT67), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT67), .B1(new_n377), .B2(new_n383), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  INV_X1    g194(.A(new_n318), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n377), .B(new_n383), .C1(new_n312), .C2(new_n313), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(KEYINPUT4), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n398), .A3(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n390), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n395), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n387), .A3(new_n389), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n384), .B(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n408), .B2(new_n396), .ZN(new_n409));
  INV_X1    g208(.A(new_n389), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n388), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n364), .B(new_n370), .C1(new_n403), .C2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n401), .A2(new_n402), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n414), .A2(new_n390), .B1(new_n406), .B2(new_n411), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n415), .B2(new_n370), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n369), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n413), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G8gat), .B(G36gat), .Z(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT64), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT24), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(G183gat), .A3(G190gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G183gat), .B(G190gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n423), .B(new_n425), .C1(new_n426), .C2(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n424), .ZN(new_n429));
  INV_X1    g228(.A(G169gat), .ZN(new_n430));
  INV_X1    g229(.A(G176gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT23), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT23), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(G169gat), .B2(G176gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n425), .ZN(new_n438));
  INV_X1    g237(.A(G183gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G190gat), .ZN(new_n440));
  INV_X1    g239(.A(G190gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G183gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n443), .B2(KEYINPUT24), .ZN(new_n444));
  INV_X1    g243(.A(new_n436), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n444), .B(new_n445), .C1(new_n423), .C2(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n435), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n431), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(KEYINPUT26), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n449), .A2(KEYINPUT26), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n450), .A2(new_n451), .B1(G183gat), .B2(G190gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(KEYINPUT27), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT27), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G183gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n441), .A2(KEYINPUT28), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(G190gat), .B1(new_n453), .B2(KEYINPUT65), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT28), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n452), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n315), .ZN(new_n468));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(KEYINPUT73), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n294), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n467), .B2(new_n315), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n447), .B2(new_n466), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n334), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n422), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n476), .A3(new_n422), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT30), .A4(new_n422), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n419), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n394), .A2(new_n467), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n393), .A2(new_n447), .A3(new_n466), .ZN(new_n487));
  INV_X1    g286(.A(G227gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(new_n278), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G71gat), .B(G99gat), .Z(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT33), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(KEYINPUT32), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n486), .A2(new_n487), .A3(new_n489), .A4(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(KEYINPUT32), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n487), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n489), .A2(KEYINPUT34), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  AOI211_X1 g307(.A(KEYINPUT70), .B(new_n508), .C1(new_n486), .C2(new_n487), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n393), .A2(new_n447), .A3(new_n466), .ZN(new_n511));
  INV_X1    g310(.A(new_n391), .ZN(new_n512));
  INV_X1    g311(.A(new_n392), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n447), .A2(new_n466), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT69), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n486), .A2(new_n516), .A3(new_n487), .ZN(new_n517));
  INV_X1    g316(.A(new_n489), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT34), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n495), .B1(new_n499), .B2(new_n494), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n490), .A2(KEYINPUT32), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n497), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n520), .A3(new_n510), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n521), .A3(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n363), .A2(new_n485), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT88), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n363), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n369), .B(KEYINPUT85), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n417), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n416), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n369), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(KEYINPUT87), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(KEYINPUT87), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n522), .A2(new_n526), .ZN(new_n545));
  INV_X1    g344(.A(new_n484), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n537), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n536), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n414), .A2(new_n387), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n410), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n409), .A2(new_n410), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT39), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n538), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n554), .B(new_n555), .C1(KEYINPUT39), .C2(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT40), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n556), .A2(new_n557), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n484), .A2(new_n539), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(KEYINPUT86), .A3(new_n557), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n477), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n422), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n566), .B1(new_n473), .B2(new_n476), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT38), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n470), .A2(new_n472), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n566), .B1(new_n572), .B2(new_n334), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n294), .B1(new_n474), .B2(new_n475), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT38), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n544), .A2(new_n479), .A3(new_n571), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n564), .A2(new_n363), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n545), .A2(KEYINPUT36), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n363), .A2(new_n485), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n275), .B1(new_n550), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n591), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n596), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n251), .A2(new_n256), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n230), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n587), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(G190gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n441), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT99), .B1(new_n607), .B2(new_n291), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(G218gat), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n589), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(new_n606), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n441), .B1(new_n601), .B2(new_n603), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n291), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND4_X1   g413(.A1(new_n611), .A2(new_n614), .A3(new_n589), .A4(new_n609), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n586), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G57gat), .B(G64gat), .Z(new_n617));
  NAND2_X1  g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT9), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n618), .A2(new_n623), .B1(new_n620), .B2(KEYINPUT98), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n379), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n240), .B1(KEYINPUT21), .B2(new_n627), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n633), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n614), .A2(new_n611), .A3(new_n609), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n588), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n608), .A2(new_n589), .A3(new_n609), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n585), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n616), .A2(new_n638), .A3(KEYINPUT101), .A4(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n627), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n600), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n598), .B1(new_n596), .B2(new_n597), .ZN(new_n652));
  INV_X1    g451(.A(new_n597), .ZN(new_n653));
  AOI211_X1 g452(.A(KEYINPUT100), .B(new_n653), .C1(new_n591), .C2(new_n595), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n627), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G120gat), .B(G148gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT103), .Z(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n647), .B1(new_n650), .B2(new_n655), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n657), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n647), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n664), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n663), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n665), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n645), .A2(new_n646), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n584), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n419), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g478(.A1(new_n676), .A2(new_n546), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n234), .B2(new_n680), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n682), .B(new_n683), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n676), .B2(new_n581), .ZN(new_n685));
  INV_X1    g484(.A(new_n545), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n676), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n363), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n536), .B2(new_n549), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n360), .A2(new_n362), .B1(new_n528), .B2(new_n529), .ZN(new_n694));
  AOI211_X1 g493(.A(KEYINPUT88), .B(new_n547), .C1(new_n694), .C2(new_n485), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n534), .B1(new_n531), .B2(KEYINPUT35), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n692), .B(new_n549), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n583), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(KEYINPUT106), .B(new_n583), .C1(new_n693), .C2(new_n698), .ZN(new_n702));
  INV_X1    g501(.A(new_n642), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n585), .B1(new_n640), .B2(new_n641), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT44), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n550), .B2(new_n583), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n638), .A2(new_n673), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n275), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n677), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n708), .A2(new_n714), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n207), .A3(new_n419), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1328gat));
  OAI21_X1  g519(.A(G36gat), .B1(new_n715), .B2(new_n546), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n208), .A3(new_n484), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n717), .A2(new_n725), .A3(new_n545), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(KEYINPUT47), .ZN(new_n727));
  INV_X1    g526(.A(new_n581), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n711), .A2(new_n728), .A3(new_n714), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730));
  OAI21_X1  g529(.A(G43gat), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n715), .A2(KEYINPUT108), .A3(new_n581), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n729), .A2(new_n725), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n726), .B(KEYINPUT107), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(G1330gat));
  OAI21_X1  g537(.A(G50gat), .B1(new_n715), .B2(new_n363), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT110), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n363), .A2(G50gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n713), .A2(new_n705), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n584), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n711), .A2(new_n537), .A3(new_n714), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n355), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n740), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n739), .B(new_n745), .C1(KEYINPUT110), .C2(KEYINPUT48), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n701), .A2(new_n702), .ZN(new_n752));
  AND4_X1   g551(.A1(new_n275), .A2(new_n645), .A3(new_n646), .A4(new_n673), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n419), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n753), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n546), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n754), .A2(new_n763), .A3(new_n545), .ZN(new_n764));
  OAI21_X1  g563(.A(G71gat), .B1(new_n757), .B2(new_n581), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n757), .A2(new_n363), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT111), .B(G78gat), .Z(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  INV_X1    g570(.A(new_n275), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n638), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n711), .A2(new_n673), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n677), .ZN(new_n775));
  INV_X1    g574(.A(new_n699), .ZN(new_n776));
  INV_X1    g575(.A(new_n705), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n773), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT51), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n776), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n419), .A2(new_n593), .A3(new_n673), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n775), .B1(new_n783), .B2(new_n784), .ZN(G1336gat));
  INV_X1    g584(.A(new_n783), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n674), .A2(new_n546), .A3(G92gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n711), .A2(new_n484), .A3(new_n673), .A4(new_n773), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n787), .B(KEYINPUT112), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n786), .A2(new_n793), .B1(new_n789), .B2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n774), .B2(new_n581), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n686), .A2(G99gat), .A3(new_n674), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n783), .B2(new_n798), .ZN(G1338gat));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n673), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n363), .B(new_n801), .C1(new_n707), .C2(new_n710), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n363), .A2(G106gat), .A3(new_n674), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n780), .B2(new_n782), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n802), .B2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI221_X1 g608(.A(new_n806), .B1(new_n800), .B2(KEYINPUT53), .C1(new_n802), .C2(new_n803), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n275), .A2(new_n645), .A3(new_n646), .A4(new_n674), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n668), .A2(new_n815), .A3(new_n670), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n656), .A2(new_n657), .A3(new_n648), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n667), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n663), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n668), .A2(new_n815), .A3(new_n670), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n663), .A4(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n665), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n247), .B1(new_n243), .B2(new_n249), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n257), .A2(new_n241), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n824), .A2(KEYINPUT115), .B1(new_n825), .B2(new_n245), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n270), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n274), .A2(new_n273), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n275), .A2(new_n823), .B1(new_n830), .B2(new_n674), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n642), .A3(new_n616), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n823), .A2(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n703), .B2(new_n704), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n638), .B1(new_n835), .B2(KEYINPUT116), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n813), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n812), .B1(new_n839), .B2(new_n537), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n832), .A2(new_n837), .A3(new_n834), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n837), .B1(new_n832), .B2(new_n834), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(new_n638), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT117), .B(new_n363), .C1(new_n843), .C2(new_n813), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n677), .A2(new_n484), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n840), .A2(new_n545), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n363), .B1(new_n843), .B2(new_n813), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n686), .B1(new_n848), .B2(new_n812), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n845), .A4(new_n844), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n851), .A3(new_n772), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(G113gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n839), .A2(new_n677), .ZN(new_n854));
  INV_X1    g653(.A(new_n694), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n484), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n772), .A2(new_n373), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT120), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n852), .A2(G113gat), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n863), .B(new_n864), .C1(new_n859), .C2(new_n860), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  AND3_X1   g665(.A1(new_n847), .A2(new_n851), .A3(new_n673), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n673), .A2(new_n375), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n867), .A2(new_n375), .B1(new_n859), .B2(new_n868), .ZN(G1341gat));
  AND3_X1   g668(.A1(new_n847), .A2(new_n851), .A3(new_n638), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n638), .A2(new_n379), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n870), .A2(new_n379), .B1(new_n857), .B2(new_n871), .ZN(G1342gat));
  NOR3_X1   g671(.A1(new_n857), .A2(G134gat), .A3(new_n705), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT56), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n847), .A2(new_n851), .A3(new_n777), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n381), .B2(new_n875), .ZN(G1343gat));
  OR2_X1    g675(.A1(new_n854), .A2(KEYINPUT121), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n854), .A2(KEYINPUT121), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n728), .A2(new_n363), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n484), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n296), .B1(new_n882), .B2(new_n275), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n836), .A2(new_n838), .ZN(new_n884));
  INV_X1    g683(.A(new_n813), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n537), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n537), .A2(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(new_n638), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n835), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n581), .A2(new_n845), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(G141gat), .A3(new_n772), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n883), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n897), .B(new_n899), .ZN(G1344gat));
  XNOR2_X1  g699(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n889), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n363), .B1(new_n885), .B2(new_n891), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(KEYINPUT57), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n674), .A3(new_n894), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n906), .B2(new_n298), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n298), .A2(KEYINPUT59), .ZN(new_n908));
  INV_X1    g707(.A(new_n895), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n674), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n882), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n298), .A3(new_n673), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n909), .B2(new_n890), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n305), .A3(new_n638), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  AOI21_X1  g716(.A(G162gat), .B1(new_n912), .B2(new_n777), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n705), .A2(new_n306), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n895), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n546), .A2(new_n419), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n849), .A2(new_n844), .A3(new_n921), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n430), .A3(new_n275), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n839), .A2(new_n419), .A3(new_n546), .A4(new_n855), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n772), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n922), .B2(new_n674), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n431), .A3(new_n673), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n922), .B2(new_n890), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n924), .A2(new_n457), .A3(new_n459), .A4(new_n638), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n441), .A3(new_n777), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n922), .A2(new_n705), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(G190gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n938), .B2(G190gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  OR2_X1    g741(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n581), .A2(new_n921), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(new_n275), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n839), .A2(new_n419), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n880), .A2(new_n546), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n772), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n948), .A2(new_n953), .ZN(G1352gat));
  NOR3_X1   g753(.A1(new_n951), .A2(G204gat), .A3(new_n674), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n943), .A2(new_n673), .A3(new_n944), .A4(new_n945), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n957), .A2(new_n958), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(G1353gat));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n638), .ZN(new_n963));
  OAI21_X1  g762(.A(G211gat), .B1(new_n905), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  NAND3_X1  g764(.A1(new_n952), .A2(new_n331), .A3(new_n638), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(new_n291), .B1(new_n951), .B2(new_n705), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n777), .A2(G218gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n946), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n972), .B(new_n968), .C1(new_n946), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1355gat));
endmodule


