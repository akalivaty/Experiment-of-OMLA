//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1247, new_n1248;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n209), .B1(new_n213), .B2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n212), .A2(KEYINPUT65), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT66), .B(KEYINPUT0), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n218), .B(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n206), .A2(G50), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n211), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G116), .A2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G50), .ZN(new_n231));
  INV_X1    g0031(.A(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G97), .ZN(new_n233));
  INV_X1    g0033(.A(G257), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n230), .B1(new_n231), .B2(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n229), .B(new_n235), .C1(G107), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT68), .B(G244), .Z(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G77), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n212), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n225), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n220), .B(new_n241), .C1(new_n240), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n253), .B(KEYINPUT69), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G68), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G58), .B(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n223), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT71), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(G223), .B1(G77), .B2(new_n267), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n262), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT70), .B1(new_n260), .B2(new_n223), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n259), .A2(new_n276), .A3(G1), .A4(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n275), .A2(new_n277), .A3(G274), .A4(new_n281), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n211), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT72), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n289), .B1(new_n290), .B2(new_n292), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n223), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n298), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n231), .B1(new_n210), .B2(G20), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(new_n303), .B1(new_n231), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n274), .B2(new_n285), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n288), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n293), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n294), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n298), .ZN(new_n313));
  INV_X1    g0113(.A(new_n298), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n300), .ZN(new_n315));
  OAI21_X1  g0115(.A(G77), .B1(new_n211), .B2(G1), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n313), .B1(G77), .B2(new_n300), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n282), .A2(new_n237), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n284), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n272), .A2(G238), .ZN(new_n320));
  INV_X1    g0120(.A(G107), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  INV_X1    g0122(.A(G232), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n271), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n320), .B1(new_n321), .B2(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n261), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n317), .B1(new_n326), .B2(G190), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n287), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n317), .C1(G169), .C2(new_n326), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(new_n286), .B2(G190), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n286), .B2(new_n328), .ZN(new_n338));
  OAI211_X1 g0138(.A(KEYINPUT73), .B(G200), .C1(new_n274), .C2(new_n285), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n336), .A2(new_n342), .A3(new_n338), .A4(new_n339), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n308), .B(new_n332), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n281), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n275), .A2(new_n345), .A3(G232), .A4(new_n277), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G223), .A2(G1698), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n232), .B2(G1698), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n322), .B1(G33), .B2(G87), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n284), .B(new_n346), .C1(new_n349), .C2(new_n262), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G200), .B2(new_n350), .ZN(new_n353));
  INV_X1    g0153(.A(G159), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n292), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n204), .A2(new_n358), .A3(new_n205), .A4(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n264), .B2(new_n266), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n263), .A2(G33), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n211), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT16), .B(new_n361), .C1(new_n368), .C2(new_n203), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n298), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n264), .A2(new_n266), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n367), .A2(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n264), .B2(new_n371), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n264), .B2(new_n266), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n372), .A2(new_n374), .B1(new_n375), .B2(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT16), .B1(new_n377), .B2(new_n361), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT79), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n293), .B1(new_n210), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n302), .B1(new_n301), .B2(new_n293), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT80), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n362), .B1(new_n364), .B2(KEYINPUT78), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(KEYINPUT78), .B2(new_n267), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n367), .B1(new_n322), .B2(G20), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n203), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n361), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n298), .A4(new_n369), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n353), .A2(new_n379), .A3(new_n382), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n379), .A2(new_n382), .A3(new_n391), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n350), .A2(G169), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n287), .B2(new_n350), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n396), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G77), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n295), .A2(new_n409), .B1(new_n211), .B2(G68), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT74), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n291), .A2(G50), .ZN(new_n413));
  XOR2_X1   g0213(.A(new_n413), .B(KEYINPUT75), .Z(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n410), .B2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n298), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT11), .B(new_n298), .C1(new_n412), .C2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT12), .B1(new_n300), .B2(G68), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n300), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n203), .B1(new_n210), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n420), .A2(new_n421), .B1(new_n302), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n265), .A2(new_n233), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G226), .A2(G1698), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n323), .B2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(new_n322), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n428), .A2(new_n262), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n275), .A2(new_n345), .A3(G238), .A4(new_n277), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n284), .A4(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n284), .B(new_n431), .C1(new_n428), .C2(new_n262), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n351), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n328), .B1(new_n432), .B2(new_n434), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n424), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n439), .A3(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n432), .A2(new_n434), .A3(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n435), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT76), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n443), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n441), .A4(new_n440), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n438), .B1(new_n448), .B2(new_n424), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n344), .A2(new_n408), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT21), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n322), .A2(G257), .A3(new_n271), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n267), .A2(G303), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n322), .A2(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G264), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n261), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n210), .B(G45), .C1(new_n279), .C2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n279), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n278), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G270), .ZN(new_n465));
  INV_X1    g0265(.A(new_n278), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G274), .A3(new_n463), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n457), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G169), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n211), .C1(G33), .C2(new_n233), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n298), .C1(new_n211), .C2(G116), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT20), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n301), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n302), .B1(G1), .B2(new_n265), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n451), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n468), .A2(G200), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n478), .C1(new_n351), .C2(new_n468), .ZN(new_n481));
  AND4_X1   g0281(.A1(G179), .A2(new_n457), .A3(new_n465), .A4(new_n467), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n473), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(KEYINPUT21), .A3(new_n468), .A4(G169), .ZN(new_n485));
  AND4_X1   g0285(.A1(new_n479), .A2(new_n481), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n322), .A2(G250), .A3(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n322), .A2(G244), .A3(new_n271), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n470), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT4), .B1(new_n268), .B2(G244), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n261), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n464), .A2(G257), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n467), .A3(new_n493), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n321), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n233), .A2(new_n321), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n376), .A2(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n314), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n301), .A2(new_n233), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n476), .B2(new_n233), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n494), .A2(new_n306), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n495), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n227), .A2(KEYINPUT85), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n322), .A2(new_n211), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n321), .A3(G20), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n516), .C1(new_n474), .C2(new_n294), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT86), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n513), .A2(new_n518), .A3(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n511), .B(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT86), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n517), .B(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n298), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n278), .A2(new_n463), .A3(new_n455), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n322), .A2(G257), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT89), .B(G294), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n528), .A2(new_n271), .B1(new_n265), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT88), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n324), .B2(new_n228), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n322), .A2(KEYINPUT88), .A3(G250), .A4(new_n271), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n467), .B(new_n527), .C1(new_n534), .C2(new_n262), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n533), .ZN(new_n537));
  INV_X1    g0337(.A(new_n530), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n261), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(G190), .A3(new_n467), .A4(new_n527), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT87), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT25), .ZN(new_n543));
  AOI211_X1 g0343(.A(G107), .B(new_n300), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  INV_X1    g0347(.A(new_n476), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n547), .B1(G107), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n525), .A2(new_n536), .A3(new_n541), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n494), .A2(G200), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n506), .C1(new_n351), .C2(new_n494), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n509), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n322), .A2(G238), .A3(new_n271), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(G244), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n454), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n261), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n210), .A2(G45), .ZN(new_n559));
  MUX2_X1   g0359(.A(G274), .B(G250), .S(new_n559), .Z(new_n560));
  NAND2_X1  g0360(.A1(new_n466), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G200), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n311), .A2(new_n301), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n294), .B2(new_n233), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n322), .A2(new_n211), .ZN(new_n568));
  NOR3_X1   g0368(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT83), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(new_n425), .B2(KEYINPUT19), .ZN(new_n571));
  OAI221_X1 g0371(.A(new_n567), .B1(new_n203), .B2(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n565), .B1(new_n572), .B2(new_n298), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n548), .A2(G87), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n557), .A2(new_n261), .B1(new_n466), .B2(new_n560), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n563), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n570), .A2(new_n571), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n567), .B1(new_n568), .B2(new_n203), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n298), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n311), .B(KEYINPUT84), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(new_n476), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n582), .A3(new_n564), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n562), .A2(new_n306), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n575), .A2(new_n287), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n526), .B1(new_n539), .B2(new_n261), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n287), .A3(new_n467), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n535), .A2(new_n306), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT24), .B1(new_n513), .B2(new_n518), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n521), .A2(new_n523), .A3(new_n520), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n314), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n549), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n589), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n553), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n450), .A2(new_n486), .A3(new_n597), .ZN(G372));
  AND3_X1   g0398(.A1(new_n509), .A2(new_n550), .A3(new_n552), .ZN(new_n599));
  INV_X1    g0399(.A(new_n586), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n573), .A2(new_n574), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT91), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n573), .A2(new_n603), .A3(new_n574), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n563), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n562), .A2(KEYINPUT90), .A3(G200), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(new_n576), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n600), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n485), .A2(new_n484), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n479), .ZN(new_n612));
  INV_X1    g0412(.A(new_n595), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n599), .B(new_n610), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n509), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n587), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT26), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n614), .A2(new_n586), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n450), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n438), .A2(new_n331), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n448), .B2(new_n424), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n399), .A2(new_n406), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n405), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n341), .A2(new_n343), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n308), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(G369));
  NAND3_X1  g0428(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT92), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G343), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n483), .ZN(new_n637));
  MUX2_X1   g0437(.A(new_n612), .B(new_n486), .S(new_n637), .Z(new_n638));
  INV_X1    g0438(.A(KEYINPUT93), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n593), .A2(new_n594), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n550), .B1(new_n643), .B2(new_n635), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n595), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n613), .A2(new_n635), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n612), .A2(new_n635), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT94), .Z(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n646), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n217), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n570), .A2(new_n474), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n210), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n221), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g0459(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n620), .A2(new_n635), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(KEYINPUT29), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n482), .A2(new_n588), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n575), .A2(new_n492), .A3(new_n467), .A4(new_n493), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n666), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(KEYINPUT30), .A3(new_n482), .A4(new_n588), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n575), .A2(G179), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n535), .A2(new_n670), .A3(new_n494), .A4(new_n468), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n636), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT31), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n636), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n587), .A2(new_n595), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n599), .A2(new_n678), .A3(new_n486), .A4(new_n635), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT96), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n597), .A2(new_n681), .A3(new_n486), .A4(new_n635), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n610), .A2(new_n615), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n615), .A2(new_n618), .A3(new_n587), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n614), .A2(new_n688), .A3(new_n586), .A4(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n686), .B1(new_n690), .B2(new_n635), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n663), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n661), .B1(new_n692), .B2(G1), .ZN(G364));
  XNOR2_X1  g0493(.A(new_n641), .B(KEYINPUT98), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n656), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n215), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n210), .B1(new_n697), .B2(G45), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n640), .A2(G330), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT97), .Z(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n215), .A2(new_n265), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT100), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n638), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n655), .A2(new_n474), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT99), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n267), .B1(new_n710), .B2(G355), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n710), .B2(G355), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n655), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n222), .A2(new_n280), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n217), .A2(new_n267), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n257), .B2(G45), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n223), .B1(G20), .B2(new_n306), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n706), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n699), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR4_X1   g0521(.A1(new_n211), .A2(new_n328), .A3(G179), .A4(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n321), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT102), .B(G159), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G179), .A2(G200), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(G20), .A3(new_n351), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n211), .B1(new_n726), .B2(G190), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(KEYINPUT32), .B1(new_n233), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G190), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n724), .B(new_n731), .C1(G68), .C2(new_n733), .ZN(new_n734));
  NOR4_X1   g0534(.A1(new_n211), .A2(new_n287), .A3(new_n351), .A4(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n322), .B1(new_n736), .B2(new_n202), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n211), .A2(new_n351), .A3(new_n328), .A4(G179), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n732), .A2(new_n351), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n739), .A2(new_n227), .B1(new_n231), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n737), .B(new_n742), .C1(KEYINPUT32), .C2(new_n729), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n211), .A2(new_n287), .A3(G190), .A4(G200), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n734), .B(new_n743), .C1(new_n409), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n744), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  INV_X1    g0550(.A(G329), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n727), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n322), .B(new_n752), .C1(G322), .C2(new_n735), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n733), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n730), .ZN(new_n758));
  INV_X1    g0558(.A(new_n529), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n738), .A2(G303), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n722), .A2(G283), .B1(G326), .B2(new_n740), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n753), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n748), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n721), .B1(new_n763), .B2(new_n718), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n700), .A2(new_n703), .B1(new_n708), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n636), .A2(new_n317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n329), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n331), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n331), .A2(new_n636), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n662), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n620), .A2(new_n773), .A3(new_n635), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n699), .B1(new_n776), .B2(new_n685), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n680), .A2(new_n682), .ZN(new_n778));
  INV_X1    g0578(.A(new_n677), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G330), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n777), .A2(KEYINPUT105), .B1(new_n781), .B2(new_n775), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(KEYINPUT105), .B2(new_n777), .ZN(new_n783));
  INV_X1    g0583(.A(new_n718), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n704), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n699), .B1(G77), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n733), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n290), .ZN(new_n788));
  INV_X1    g0588(.A(G143), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n736), .A2(new_n789), .B1(new_n790), .B2(new_n741), .ZN(new_n791));
  INV_X1    g0591(.A(new_n725), .ZN(new_n792));
  INV_X1    g0592(.A(new_n747), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n788), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n723), .A2(new_n203), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n322), .B1(new_n798), .B2(new_n727), .C1(new_n739), .C2(new_n231), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(G58), .C2(new_n758), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n723), .A2(new_n227), .B1(new_n750), .B2(new_n727), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT104), .Z(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n739), .A2(new_n321), .B1(new_n804), .B2(new_n741), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT103), .B(G283), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n733), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n267), .B1(new_n730), .B2(new_n233), .C1(new_n736), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n793), .B2(G116), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n803), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n786), .B1(new_n813), .B2(new_n718), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n773), .B2(new_n705), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n783), .A2(new_n815), .ZN(G384));
  OR2_X1    g0616(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n817), .A2(G116), .A3(new_n224), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  NAND4_X1  g0620(.A1(new_n221), .A2(G77), .A3(new_n358), .A4(new_n359), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n231), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n210), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n400), .A2(new_n634), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT107), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n400), .A2(KEYINPUT107), .A3(new_n634), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n392), .B(KEYINPUT17), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n405), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n400), .A2(KEYINPUT107), .A3(new_n634), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT107), .B1(new_n400), .B2(new_n634), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n403), .A2(new_n392), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n829), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT108), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n836), .A2(KEYINPUT108), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT38), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n361), .B1(new_n368), .B2(new_n203), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT106), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT16), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n370), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n381), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n634), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n407), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n402), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n855), .B2(new_n852), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n856), .B2(new_n393), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n839), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT109), .B1(new_n844), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n424), .A2(new_n636), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n444), .B2(new_n447), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n449), .B2(new_n861), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NOR4_X1   g0664(.A1(new_n683), .A2(new_n863), .A3(new_n864), .A4(new_n771), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n834), .A2(KEYINPUT37), .A3(new_n835), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n837), .B1(new_n829), .B2(new_n838), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n841), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n831), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n843), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT109), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n860), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n683), .A2(new_n771), .A3(new_n863), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n854), .B2(new_n858), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n859), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n864), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n450), .A2(new_n780), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(G330), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n844), .B2(new_n859), .ZN(new_n887));
  INV_X1    g0687(.A(new_n878), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n448), .A2(new_n424), .A3(new_n635), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n405), .A2(new_n634), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n874), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n863), .B1(new_n774), .B2(new_n770), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n450), .B1(new_n663), .B2(new_n691), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n627), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n885), .A2(new_n899), .B1(new_n210), .B2(new_n697), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT110), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n885), .A2(new_n899), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n824), .B1(new_n902), .B2(new_n904), .ZN(G367));
  NAND3_X1  g0705(.A1(new_n636), .A2(new_n602), .A3(new_n604), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n610), .A2(KEYINPUT111), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n586), .B2(new_n906), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT111), .B1(new_n610), .B2(new_n906), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n706), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n719), .B1(new_n217), .B2(new_n311), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n715), .A2(new_n249), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n699), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n793), .A2(new_n807), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n267), .B1(new_n736), .B2(new_n804), .ZN(new_n916));
  INV_X1    g0716(.A(new_n727), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(G317), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n723), .A2(new_n233), .B1(new_n529), .B2(new_n787), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n741), .A2(new_n750), .B1(new_n730), .B2(new_n321), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n738), .A2(G116), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n915), .A2(new_n918), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n793), .A2(G50), .B1(new_n792), .B2(new_n733), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT115), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n322), .B1(new_n727), .B2(new_n790), .C1(new_n736), .C2(new_n290), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n739), .A2(new_n202), .B1(new_n723), .B2(new_n409), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n741), .A2(new_n789), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n730), .A2(new_n203), .ZN(new_n930));
  NOR4_X1   g0730(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n925), .A2(KEYINPUT115), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT47), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n914), .B1(new_n935), .B2(new_n718), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n911), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n698), .B(KEYINPUT114), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT113), .B1(new_n650), .B2(new_n647), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(new_n651), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(new_n641), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n694), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n509), .A2(new_n635), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT112), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n509), .B(new_n552), .C1(new_n506), .C2(new_n635), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n652), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n653), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n652), .B2(new_n950), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n648), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n953), .A2(new_n957), .A3(new_n648), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n945), .A2(new_n960), .A3(new_n692), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n692), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n656), .B(KEYINPUT41), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n939), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n509), .B1(new_n950), .B2(new_n595), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n650), .A2(new_n647), .A3(new_n949), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n967), .A2(new_n635), .B1(new_n968), .B2(KEYINPUT42), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n910), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n969), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n972), .B(new_n973), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n648), .A2(new_n950), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n937), .B1(new_n966), .B2(new_n977), .ZN(G387));
  NOR3_X1   g0778(.A1(new_n246), .A2(new_n280), .A3(new_n322), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n293), .B2(G50), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n309), .A2(new_n980), .A3(new_n231), .ZN(new_n983));
  AOI21_X1  g0783(.A(G45), .B1(G68), .B2(G77), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n657), .B1(new_n985), .B2(new_n267), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n217), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n719), .C1(new_n321), .C2(new_n217), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n309), .A2(new_n733), .B1(G159), .B2(new_n740), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n233), .B2(new_n723), .C1(new_n409), .C2(new_n739), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n267), .B1(new_n744), .B2(G68), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n290), .B2(new_n727), .C1(new_n231), .C2(new_n736), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n581), .A2(new_n730), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n723), .A2(new_n474), .ZN(new_n995));
  INV_X1    g0795(.A(G326), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n267), .B1(new_n727), .B2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n735), .A2(G317), .B1(G311), .B2(new_n733), .ZN(new_n998));
  INV_X1    g0798(.A(G322), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n999), .B2(new_n741), .C1(new_n747), .C2(new_n804), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n738), .A2(new_n759), .B1(new_n758), .B2(new_n807), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n995), .B(new_n997), .C1(new_n1006), .C2(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n994), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n699), .B(new_n988), .C1(new_n1009), .C2(new_n784), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n647), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n706), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n945), .B2(new_n939), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n692), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n944), .A2(KEYINPUT117), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n942), .A2(new_n943), .A3(new_n692), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n656), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT117), .B1(new_n944), .B2(new_n1014), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(G393));
  INV_X1    g0819(.A(new_n961), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n648), .B1(new_n953), .B2(new_n957), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT118), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT118), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n939), .A3(new_n1024), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n253), .A2(new_n217), .A3(new_n267), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n719), .B1(new_n233), .B2(new_n217), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n699), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n735), .A2(G311), .B1(G317), .B2(new_n740), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT52), .Z(new_n1030));
  OAI21_X1  g0830(.A(new_n267), .B1(new_n727), .B2(new_n999), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G294), .B2(new_n744), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n724), .B1(G303), .B2(new_n733), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n738), .A2(new_n807), .B1(new_n758), .B2(G116), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n735), .A2(G159), .B1(G150), .B2(new_n740), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n739), .A2(new_n203), .B1(new_n231), .B2(new_n787), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n730), .A2(new_n409), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n322), .B1(new_n727), .B2(new_n789), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G87), .B2(new_n722), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n293), .C2(new_n747), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1028), .B1(new_n1044), .B2(new_n718), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n949), .B2(new_n707), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n962), .A2(new_n1047), .A3(new_n656), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1025), .A2(new_n1046), .A3(new_n1048), .ZN(G390));
  NOR3_X1   g0849(.A1(new_n781), .A2(new_n771), .A3(new_n863), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n690), .A2(new_n635), .A3(new_n769), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n770), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n863), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n890), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n860), .A2(new_n875), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n894), .A2(new_n890), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n887), .B2(new_n889), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1050), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n860), .A2(new_n875), .A3(new_n1054), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n683), .A2(new_n684), .A3(new_n771), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n1053), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT39), .B1(new_n872), .B2(new_n874), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n859), .A2(new_n878), .A3(new_n886), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1059), .B(new_n1061), .C1(new_n1064), .C2(new_n1056), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n450), .A2(new_n685), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n897), .A2(new_n627), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT119), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n863), .C1(new_n781), .C2(new_n771), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT119), .B1(new_n1060), .B2(new_n1053), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1052), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1061), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n774), .A2(new_n770), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1060), .A2(new_n1053), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1050), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1068), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1066), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1058), .A2(new_n1065), .A3(new_n1077), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n656), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1058), .A2(new_n1065), .A3(new_n939), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n699), .B1(new_n309), .B2(new_n785), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n267), .B1(new_n727), .B2(new_n809), .C1(new_n736), .C2(new_n474), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n797), .B(new_n1084), .C1(G87), .C2(new_n738), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n233), .B2(new_n747), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1039), .B1(new_n733), .B2(G107), .ZN(new_n1087));
  INV_X1    g0887(.A(G283), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n741), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT120), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n322), .B1(new_n727), .B2(new_n1092), .C1(new_n736), .C2(new_n798), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n793), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n738), .A2(G150), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT53), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n758), .A2(G159), .B1(G137), .B2(new_n733), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n722), .A2(G50), .B1(G128), .B2(new_n740), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1090), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1083), .B1(new_n1103), .B2(new_n718), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1064), .B2(new_n705), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1082), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1081), .A2(new_n1106), .ZN(G378));
  OAI21_X1  g0907(.A(new_n699), .B1(G50), .B2(new_n785), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n305), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(new_n852), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n308), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n626), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n308), .B(new_n1110), .C1(new_n341), .C2(new_n343), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n705), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n322), .A2(G41), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G50), .B(new_n1121), .C1(new_n265), .C2(new_n279), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n1088), .B2(new_n727), .C1(new_n736), .C2(new_n321), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n930), .B(new_n1123), .C1(G77), .C2(new_n738), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n723), .A2(new_n202), .B1(new_n474), .B2(new_n741), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G97), .B2(new_n733), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(new_n581), .C2(new_n749), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT58), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n749), .A2(new_n790), .B1(new_n1092), .B2(new_n741), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n787), .A2(new_n798), .B1(new_n730), .B2(new_n290), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G128), .A2(new_n735), .B1(new_n738), .B2(new_n1095), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1130), .B(new_n1131), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT59), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G33), .B(G41), .C1(new_n917), .C2(G124), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n725), .B2(new_n723), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1108), .B(new_n1120), .C1(new_n718), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n684), .B1(new_n879), .B2(new_n864), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n876), .A2(new_n1142), .A3(new_n1119), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1119), .B1(new_n876), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n896), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n876), .A2(new_n1142), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1119), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n896), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n876), .A2(new_n1142), .A3(new_n1119), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1141), .B1(new_n1152), .B2(new_n939), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1068), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1080), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n1155), .A3(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n656), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(G375));
  AND2_X1   g0959(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n938), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n863), .A2(new_n215), .A3(new_n265), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n699), .B1(G68), .B2(new_n785), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n739), .A2(new_n233), .B1(new_n809), .B2(new_n741), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n723), .A2(new_n409), .B1(new_n474), .B2(new_n787), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n747), .A2(new_n321), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n267), .B1(new_n727), .B2(new_n804), .C1(new_n736), .C2(new_n1088), .ZN(new_n1168));
  OR4_X1    g0968(.A1(new_n993), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n739), .A2(new_n354), .B1(new_n231), .B2(new_n730), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G132), .B2(new_n740), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n267), .B1(new_n917), .B2(G128), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n735), .A2(G137), .B1(new_n744), .B2(G150), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n733), .A2(new_n1095), .B1(new_n722), .B2(G58), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1163), .B1(new_n1176), .B2(new_n718), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1161), .B1(new_n1162), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1160), .A2(new_n1068), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n965), .A3(new_n1078), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(G381));
  OAI211_X1 g0981(.A(new_n765), .B(new_n1013), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1182));
  OR3_X1    g0982(.A1(G390), .A2(G384), .A3(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(G375), .A2(G378), .ZN(new_n1184));
  OR4_X1    g0984(.A1(G387), .A2(new_n1183), .A3(new_n1184), .A4(G381), .ZN(G407));
  INV_X1    g0985(.A(G343), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(G213), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT122), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g0990(.A(G390), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT125), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(G393), .A2(G396), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G387), .A2(new_n1192), .B1(new_n1182), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1014), .B1(new_n1022), .B2(new_n945), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n938), .B1(new_n1195), .B2(new_n964), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1196), .A2(new_n976), .B1(new_n911), .B2(new_n936), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1182), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1197), .B2(KEYINPUT125), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(G387), .A2(new_n1182), .A3(new_n1193), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(G390), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT61), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1186), .A2(G213), .A3(G2897), .ZN(new_n1206));
  INV_X1    g1006(.A(G384), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1160), .A2(KEYINPUT60), .A3(new_n1068), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n656), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1179), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1178), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1210), .A2(new_n1179), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G384), .B(new_n1178), .C1(new_n1214), .C2(new_n1209), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1213), .A2(KEYINPUT124), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT124), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1206), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1206), .B2(new_n1216), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G375), .A2(G378), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1152), .A2(new_n1155), .A3(new_n965), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1153), .A2(new_n1221), .A3(new_n1081), .A4(new_n1106), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n1187), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1204), .B(new_n1205), .C1(new_n1219), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1220), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT123), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT123), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1220), .A2(new_n1223), .A3(new_n1226), .A4(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n1225), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1205), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1228), .A2(new_n1236), .A3(new_n1237), .A4(new_n1231), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1224), .A2(KEYINPUT62), .A3(new_n1226), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1228), .A2(new_n1237), .A3(new_n1231), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT126), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1235), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT127), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1204), .B(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1234), .B1(new_n1243), .B2(new_n1245), .ZN(G405));
  NAND2_X1  g1046(.A1(new_n1184), .A2(new_n1220), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(new_n1226), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1245), .B(new_n1248), .ZN(G402));
endmodule


