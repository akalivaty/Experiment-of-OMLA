//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n469), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n472), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n469), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n482), .B(new_n485), .C1(G124), .C2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n464), .A2(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n469), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n505), .A2(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n503), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(G51), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n508), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(G168));
  AOI22_X1  g098(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n502), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n505), .A2(new_n526), .B1(new_n511), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  AOI22_X1  g104(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n502), .ZN(new_n531));
  INV_X1    g106(.A(G43), .ZN(new_n532));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n505), .A2(new_n532), .B1(new_n511), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  NAND3_X1  g115(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT9), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT9), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n504), .A2(new_n543), .A3(G53), .A4(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n511), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT71), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(G91), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(G65), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n519), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  OR2_X1    g129(.A1(KEYINPUT72), .A2(G65), .ZN(new_n555));
  NAND2_X1  g130(.A1(KEYINPUT72), .A2(G65), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n500), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n550), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n545), .B(new_n549), .C1(new_n554), .C2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n502), .B1(new_n519), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n505), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n547), .A2(G87), .A3(new_n548), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  OAI21_X1  g148(.A(G61), .B1(new_n508), .B2(new_n507), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n502), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .B1(new_n570), .B2(G48), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n547), .A2(G86), .A3(new_n548), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT76), .B(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n505), .A2(new_n581), .B1(new_n511), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n586), .A2(new_n587), .B1(new_n502), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n500), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n502), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n570), .A2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n547), .A2(G92), .A3(new_n548), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G321));
  OR2_X1    g176(.A1(G299), .A2(KEYINPUT79), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(KEYINPUT79), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(G168), .A2(new_n603), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT78), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G297));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G860), .ZN(G148));
  OAI21_X1  g186(.A(new_n603), .B1(new_n531), .B2(new_n534), .ZN(new_n612));
  INV_X1    g187(.A(new_n599), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n614), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n496), .A2(new_n473), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n486), .A2(G123), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n480), .A2(G135), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n622), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n638), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n649), .A2(new_n645), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n632), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n641), .A2(new_n646), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(new_n631), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n654), .A3(G14), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n686), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n687), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT26), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G129), .B2(new_n486), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n698), .A2(new_n699), .B1(new_n480), .B2(G141), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G32), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT83), .B(G29), .Z(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G34), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n478), .B2(new_n707), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n711), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(G171), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G5), .B2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n720), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT93), .B(G1966), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n713), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G27), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n729), .B(new_n734), .C1(new_n727), .C2(new_n728), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n730), .A2(G35), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n730), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n707), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n480), .A2(G139), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n496), .A2(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n469), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(new_n707), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2072), .Z(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n751), .B(new_n757), .C1(new_n627), .C2(new_n713), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n719), .A2(new_n735), .A3(new_n740), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G299), .A2(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n720), .A2(G20), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT23), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT96), .B(G1956), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n722), .A2(new_n723), .B1(new_n712), .B2(new_n718), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n709), .B2(new_n710), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT94), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n759), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n713), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT88), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G128), .B2(new_n486), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n480), .A2(G140), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT87), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2067), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n599), .B2(G16), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G1348), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(G1348), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n720), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n535), .B2(new_n720), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  NAND4_X1  g363(.A1(new_n781), .A2(new_n784), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT90), .Z(new_n790));
  NAND2_X1  g365(.A1(G288), .A2(KEYINPUT85), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT85), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n571), .A2(new_n572), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n720), .A2(G23), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT86), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT86), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n720), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n720), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1971), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n804), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n800), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n800), .A2(new_n812), .A3(new_n801), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n486), .A2(G119), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT84), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G107), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G131), .B2(new_n480), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G25), .B(new_n820), .S(new_n730), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  OR2_X1    g398(.A1(G16), .A2(G24), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G290), .B2(new_n720), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n811), .A2(new_n813), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n769), .B(new_n790), .C1(new_n831), .C2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n769), .A2(new_n790), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  AOI22_X1  g411(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n502), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n500), .A2(new_n504), .A3(G93), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n839), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n535), .B1(new_n844), .B2(KEYINPUT98), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(KEYINPUT98), .B2(new_n844), .ZN(new_n849));
  INV_X1    g424(.A(new_n844), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n535), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n599), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n847), .B1(new_n861), .B2(new_n862), .ZN(G145));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n776), .A2(new_n864), .A3(new_n778), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n776), .B2(new_n778), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(new_n748), .B2(new_n745), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n749), .A3(new_n865), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n820), .B(new_n618), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(G126), .A2(G2105), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n464), .B2(new_n465), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n469), .A2(G114), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT101), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n488), .A2(new_n881), .A3(new_n492), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n497), .B1(new_n480), .B2(G138), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n880), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n706), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n705), .A2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n486), .A2(G130), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n469), .A2(KEYINPUT103), .A3(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT103), .B1(new_n469), .B2(G118), .ZN(new_n891));
  OR2_X1    g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n890), .A2(G2104), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n480), .A2(G142), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n887), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n887), .B2(new_n888), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n873), .A2(new_n874), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n868), .A2(new_n870), .ZN(new_n901));
  INV_X1    g476(.A(new_n871), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n897), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n898), .A4(new_n872), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n627), .B(new_n478), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(G162), .Z(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n900), .A2(new_n905), .ZN(new_n911));
  INV_X1    g486(.A(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n559), .A2(new_n560), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n917), .A2(new_n561), .A3(new_n599), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n599), .B1(new_n917), .B2(new_n561), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n613), .B1(new_n562), .B2(new_n563), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n561), .A3(new_n599), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n853), .B(new_n614), .Z(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G303), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n794), .B(G305), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n927), .B(new_n929), .C1(new_n937), .C2(new_n938), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n931), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n931), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n844), .A2(new_n603), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  AOI21_X1  g521(.A(G168), .B1(G301), .B2(KEYINPUT105), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(KEYINPUT105), .B2(G301), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  NAND3_X1  g524(.A1(G171), .A2(G168), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n853), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n849), .A3(new_n852), .A4(new_n950), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n928), .A3(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n920), .A2(new_n923), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n953), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n924), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n936), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(new_n954), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n932), .B(new_n933), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n936), .B1(new_n955), .B2(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n965), .A3(new_n954), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n909), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n963), .B1(new_n959), .B2(KEYINPUT106), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n955), .A2(new_n956), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n969), .A2(new_n909), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n961), .A2(new_n979), .A3(new_n966), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n966), .A2(new_n962), .A3(new_n968), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n973), .B1(new_n983), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n885), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT109), .B(G40), .Z(new_n989));
  OAI211_X1 g564(.A(new_n468), .B(new_n989), .C1(new_n476), .C2(new_n477), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2067), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n779), .B(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n705), .B(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n820), .B(new_n822), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(G290), .B(G1986), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT113), .B(G8), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n990), .A2(G2084), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT50), .B1(new_n885), .B2(new_n985), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G164), .A2(new_n1004), .A3(G1384), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1002), .B(KEYINPUT116), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n990), .B1(new_n986), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n495), .A2(new_n498), .ZN(new_n1013));
  INV_X1    g588(.A(new_n493), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(new_n987), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n985), .A4(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n985), .A3(new_n1017), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT115), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1966), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1001), .B1(new_n1010), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n1024), .B2(G168), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1008), .A2(new_n1009), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NOR4_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(G286), .A4(new_n1001), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n990), .A2(G2090), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT111), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1034));
  INV_X1    g609(.A(new_n990), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT110), .B(G1971), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1031), .B(new_n1040), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1033), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G166), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1048), .B2(KEYINPUT55), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1030), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1042), .A2(G8), .A3(new_n1050), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n791), .A2(G1976), .A3(new_n793), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1001), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n986), .B2(new_n990), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT52), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n885), .A2(new_n985), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1001), .B1(new_n1058), .B2(new_n1035), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1059), .B(new_n1061), .C1(new_n1060), .C2(new_n794), .ZN(new_n1062));
  INV_X1    g637(.A(G1981), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n577), .A2(new_n578), .A3(new_n1063), .A4(new_n579), .ZN(new_n1064));
  INV_X1    g639(.A(G48), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT114), .B(G86), .Z(new_n1066));
  OAI22_X1  g641(.A1(new_n505), .A2(new_n1065), .B1(new_n511), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G1981), .B1(new_n1067), .B2(new_n576), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1059), .A3(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1057), .A2(new_n1062), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1052), .A2(new_n1053), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n1029), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1004), .B1(new_n885), .B2(new_n985), .ZN(new_n1077));
  NOR3_X1   g652(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n990), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1079), .A2(new_n1080), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1051), .B1(new_n1081), .B2(new_n1001), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1074), .A2(new_n1053), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1030), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1074), .A2(new_n1053), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1032), .A2(KEYINPUT111), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1044), .B1(new_n1087), .B2(new_n1041), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT63), .B1(new_n1088), .B2(new_n1050), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n1091), .C1(new_n1028), .C2(new_n1025), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1076), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1073), .A2(new_n1060), .A3(new_n572), .A4(new_n571), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1056), .B1(new_n1094), .B2(new_n1064), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1053), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1074), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n559), .B(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1956), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1015), .A2(new_n1004), .A3(new_n985), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1035), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(new_n1077), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n986), .A2(G2067), .A3(new_n990), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1035), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n613), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n1099), .A3(new_n1105), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1106), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1078), .A2(new_n990), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1077), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1956), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n559), .B(KEYINPUT57), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n1035), .A2(new_n1034), .A3(new_n1036), .A4(new_n1104), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1114), .B1(new_n1120), .B2(new_n1106), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n986), .B2(new_n990), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1037), .B2(G1996), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n535), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1129), .A3(new_n535), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1128), .A2(new_n1130), .B1(new_n1110), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1110), .A2(new_n613), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1133), .B2(new_n1111), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT119), .B(new_n1114), .C1(new_n1120), .C2(new_n1106), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1118), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1112), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1113), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1037), .B2(G2078), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1108), .A2(new_n723), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n733), .A2(KEYINPUT53), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1144), .C1(new_n1021), .C2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n1146), .B2(G171), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT123), .B(G2078), .Z(new_n1149));
  AND3_X1   g724(.A1(new_n1149), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n988), .A2(G160), .A3(new_n1034), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(G301), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1148), .A2(G301), .A3(new_n1151), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1146), .A2(G171), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1074), .A2(new_n1053), .A3(new_n1082), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1153), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1141), .A2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1026), .A2(G168), .A3(new_n1001), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G168), .A2(new_n1001), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1162), .A2(KEYINPUT51), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1024), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1044), .B1(new_n1010), .B2(new_n1023), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT51), .B1(new_n1165), .B2(new_n1162), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1166), .B2(KEYINPUT121), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(KEYINPUT51), .C1(new_n1165), .C2(new_n1162), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1161), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1093), .B(new_n1097), .C1(new_n1160), .C2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1158), .A2(new_n1156), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g749(.A(KEYINPUT62), .B(new_n1161), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1000), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n991), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n996), .A2(new_n822), .A3(new_n815), .A4(new_n819), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n776), .A2(new_n992), .A3(new_n778), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT124), .Z(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT46), .B1(new_n991), .B2(new_n994), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT125), .Z(new_n1184));
  NAND3_X1  g759(.A1(new_n991), .A2(KEYINPUT46), .A3(new_n994), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT126), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1178), .B1(new_n993), .B2(new_n706), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1178), .A2(G1986), .A3(G290), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT48), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n991), .B2(new_n998), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1182), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1177), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n461), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n655), .B(new_n1197), .C1(new_n691), .C2(new_n692), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1198), .B1(new_n910), .B2(new_n913), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n972), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1196), .B1(new_n972), .B2(new_n1199), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n1201), .ZN(G308));
  NAND2_X1  g776(.A1(new_n972), .A2(new_n1199), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(KEYINPUT127), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n972), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(G225));
endmodule


