//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n469), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n469), .A2(new_n476), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n465), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G102), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n476), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT3), .B(G2104), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G138), .A4(new_n476), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n497), .A2(new_n499), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n512), .A2(new_n513), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n507), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(new_n511), .B1(new_n528), .B2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n515), .A2(new_n534), .B1(new_n517), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n511), .A2(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n521), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n540));
  OR3_X1    g115(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n536), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n515), .A2(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(new_n511), .A2(G65), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT71), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n515), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G91), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n528), .A2(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g142(.A(new_n562), .B(new_n563), .C1(new_n528), .C2(G53), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n559), .B(new_n561), .C1(new_n567), .C2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  OR2_X1    g145(.A1(new_n519), .A2(new_n522), .ZN(G303));
  NAND2_X1  g146(.A1(new_n560), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n528), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n511), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT72), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n521), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G86), .B2(new_n560), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n528), .A2(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n528), .A2(G47), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT73), .B(G85), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n515), .B2(new_n584), .C1(new_n585), .C2(new_n521), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT10), .B1(new_n515), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n508), .A2(new_n510), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n596), .B(KEYINPUT74), .C1(new_n597), .C2(new_n517), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n517), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n591), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n587), .B1(G868), .B2(new_n602), .ZN(G284));
  OAI21_X1  g178(.A(new_n587), .B1(G868), .B2(new_n602), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT75), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT76), .Z(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n503), .A2(new_n498), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2100), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n484), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n480), .A2(G135), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2435), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2438), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  AOI21_X1  g227(.A(KEYINPUT18), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n650), .B(new_n653), .Z(G227));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT77), .ZN(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n656), .A2(new_n657), .ZN(new_n663));
  AOI22_X1  g238(.A1(new_n661), .A2(new_n662), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n658), .A2(new_n663), .A3(new_n660), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(new_n662), .C2(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G21), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n674), .A2(G16), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G286), .B2(G16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT90), .ZN(new_n677));
  INV_X1    g252(.A(G1966), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G35), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G162), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT29), .Z(new_n683));
  INV_X1    g258(.A(G2090), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT93), .ZN(new_n686));
  MUX2_X1   g261(.A(G22), .B(G303), .S(G16), .Z(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G23), .B(G288), .S(G16), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT82), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G6), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G305), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT81), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n689), .A2(new_n693), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT34), .Z(new_n701));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1986), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n680), .A2(G25), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n484), .A2(G119), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT79), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n708));
  INV_X1    g283(.A(G95), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n476), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT80), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n480), .A2(G131), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT35), .B(G1991), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n714), .A2(new_n716), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n704), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n701), .A2(new_n702), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n702), .B1(new_n701), .B2(new_n719), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n679), .B(new_n686), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(G171), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G5), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G4), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n601), .A2(new_n598), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n729), .A2(new_n590), .A3(new_n589), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1348), .ZN(new_n732));
  INV_X1    g307(.A(new_n549), .ZN(new_n733));
  MUX2_X1   g308(.A(G19), .B(new_n733), .S(G16), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n484), .A2(G128), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n480), .A2(G140), .ZN(new_n737));
  NOR2_X1   g312(.A1(G104), .A2(G2105), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n476), .B2(G116), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n680), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT83), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n732), .A2(new_n735), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT84), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n680), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G160), .B2(new_n680), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G2084), .Z(new_n755));
  NOR2_X1   g330(.A1(new_n677), .A2(new_n678), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT91), .Z(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT92), .B(G28), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(new_n680), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n626), .B2(new_n680), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n680), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT86), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G129), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n480), .A2(G141), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n498), .A2(G105), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(new_n680), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT88), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT27), .B(G1996), .Z(new_n776));
  AOI21_X1  g351(.A(new_n761), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n749), .A2(new_n755), .A3(new_n757), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n722), .A2(new_n726), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G27), .A2(G29), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2078), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT31), .B(G11), .Z(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G299), .A2(G16), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n786));
  INV_X1    g361(.A(G20), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n786), .A2(new_n787), .A3(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n683), .B2(new_n684), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT94), .Z(new_n794));
  OR2_X1    g369(.A1(new_n685), .A2(KEYINPUT93), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n779), .A2(new_n784), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n775), .A2(new_n776), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT89), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n498), .A2(G103), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n480), .A2(G139), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n476), .B2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G33), .B(new_n807), .S(G29), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2072), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n796), .A2(new_n798), .A3(new_n809), .ZN(G311));
  NOR2_X1   g385(.A1(new_n722), .A2(new_n778), .ZN(new_n811));
  INV_X1    g386(.A(new_n726), .ZN(new_n812));
  AND4_X1   g387(.A1(new_n794), .A2(new_n811), .A3(new_n795), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n798), .ZN(new_n814));
  INV_X1    g389(.A(new_n809), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n813), .A2(new_n814), .A3(new_n784), .A4(new_n815), .ZN(G150));
  XNOR2_X1  g391(.A(KEYINPUT96), .B(G860), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT95), .B(G93), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n515), .A2(new_n818), .B1(new_n517), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n521), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n817), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n820), .A2(new_n822), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n549), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n730), .A2(new_n609), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n817), .ZN(G145));
  XOR2_X1   g406(.A(KEYINPUT101), .B(G37), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n492), .B(KEYINPUT97), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n478), .ZN(new_n835));
  INV_X1    g410(.A(new_n626), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(G160), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n626), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n773), .B(new_n713), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n505), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT99), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(G164), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n807), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n484), .A2(G130), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n480), .A2(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n740), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n619), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n849), .A2(new_n855), .ZN(new_n858));
  INV_X1    g433(.A(new_n619), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n849), .A2(new_n855), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n847), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n843), .A2(new_n846), .A3(new_n857), .A4(new_n861), .ZN(new_n864));
  AOI211_X1 g439(.A(KEYINPUT100), .B(new_n840), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(new_n840), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n833), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n863), .A2(new_n840), .A3(new_n864), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT40), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n847), .A2(new_n862), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n843), .A2(new_n846), .B1(new_n857), .B2(new_n861), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n867), .A2(new_n866), .A3(new_n868), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n832), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n871), .B(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n873), .A2(new_n883), .ZN(G395));
  XOR2_X1   g459(.A(new_n549), .B(new_n825), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n613), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n602), .A2(new_n606), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n602), .A2(new_n606), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT41), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n730), .A2(G299), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n887), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n887), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n886), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(G288), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G166), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G290), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(G290), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(G305), .ZN(new_n909));
  INV_X1    g484(.A(G305), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n905), .A2(G290), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n906), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n902), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n902), .B2(new_n903), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n825), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT104), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n899), .A2(new_n921), .A3(KEYINPUT41), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n541), .A2(G168), .A3(new_n542), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G168), .B1(new_n541), .B2(new_n542), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n885), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n826), .A3(new_n924), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n924), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n931), .B2(new_n885), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n920), .B(new_n922), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n892), .A3(new_n887), .A4(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n913), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n930), .A2(new_n932), .A3(new_n899), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n909), .A2(new_n912), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n890), .A2(new_n894), .B1(new_n927), .B2(new_n929), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n942), .A3(new_n833), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT105), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n832), .B1(new_n935), .B2(new_n913), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n942), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n919), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n913), .B1(new_n937), .B2(new_n940), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(new_n919), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT44), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n951), .A2(new_n919), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n945), .B2(new_n942), .ZN(new_n956));
  OR3_X1    g531(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT44), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n953), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n954), .B1(new_n953), .B2(new_n957), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(G397));
  NAND3_X1  g535(.A1(new_n472), .A2(new_n477), .A3(G40), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  INV_X1    g537(.A(new_n495), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n503), .B2(G126), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n499), .B1(new_n964), .B2(new_n476), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n502), .A2(new_n504), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT45), .B(new_n962), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n961), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n967), .B2(new_n968), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT111), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT110), .B1(new_n969), .B2(new_n970), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  NOR4_X1   g553(.A1(new_n977), .A2(new_n978), .A3(new_n961), .A4(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n688), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n961), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n502), .A2(new_n504), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n496), .A2(G2105), .B1(G102), .B2(new_n498), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n505), .A2(new_n987), .A3(new_n962), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n684), .ZN(new_n992));
  INV_X1    g567(.A(new_n970), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n505), .B2(new_n962), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n972), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(new_n983), .A3(new_n975), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n978), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n995), .A2(KEYINPUT111), .A3(new_n975), .A4(new_n983), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT112), .A3(new_n688), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n982), .A2(new_n992), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G303), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT55), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(KEYINPUT55), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1001), .A2(G8), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n579), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G305), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(KEYINPUT115), .B2(KEYINPUT49), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n967), .A2(new_n961), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1018));
  OAI211_X1 g593(.A(new_n1014), .B(new_n1017), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(G288), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n904), .A2(G1976), .ZN(new_n1023));
  OR3_X1    g598(.A1(new_n1021), .A2(KEYINPUT52), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1020), .A3(new_n904), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(G1981), .B2(G305), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1010), .A2(new_n1026), .B1(new_n1017), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n969), .A2(new_n983), .A3(new_n970), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n678), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT118), .B(G2084), .Z(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n983), .A3(new_n989), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1016), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G286), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(KEYINPUT63), .ZN(new_n1039));
  INV_X1    g614(.A(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n997), .A2(new_n1040), .A3(new_n998), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT121), .B1(new_n988), .B2(new_n990), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1032), .A2(new_n1045), .A3(new_n983), .A4(new_n989), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n725), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT125), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT125), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1044), .A2(new_n1049), .A3(new_n725), .A4(new_n1046), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(G171), .B(KEYINPUT54), .ZN(new_n1052));
  INV_X1    g627(.A(new_n971), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n961), .B(KEYINPUT126), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT53), .A4(new_n1040), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1043), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1053), .A2(KEYINPUT53), .A3(new_n1040), .A4(new_n983), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1047), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT124), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1047), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1060), .A2(new_n1062), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1057), .B1(new_n1063), .B2(new_n1052), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G286), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT122), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n991), .A2(new_n1033), .B1(new_n678), .B2(new_n1030), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT123), .B(new_n1067), .C1(new_n1068), .C2(new_n1016), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1035), .B2(new_n1066), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1070), .B(new_n1073), .C1(new_n1035), .C2(new_n1066), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1068), .A2(new_n1067), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1064), .A2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n995), .A2(new_n983), .A3(new_n975), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n567), .B2(new_n568), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n606), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G299), .A2(new_n1082), .A3(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n987), .B1(new_n505), .B2(new_n962), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n1087), .B2(new_n961), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1032), .A2(new_n1089), .A3(new_n983), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n990), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1079), .B(new_n1086), .C1(new_n1091), .C2(G1956), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1015), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n967), .A2(new_n961), .A3(KEYINPUT120), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1095), .A2(G2067), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1044), .A2(new_n1098), .A3(new_n1046), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n602), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1086), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1956), .B1(new_n1103), .B2(new_n989), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1078), .ZN(new_n1105));
  NOR4_X1   g680(.A1(new_n977), .A2(new_n961), .A3(new_n974), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1102), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1093), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1087), .A2(KEYINPUT116), .A3(new_n961), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1089), .B1(new_n1032), .B2(new_n983), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n989), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n791), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1086), .B1(new_n1114), .B2(new_n1079), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1110), .B1(new_n1115), .B2(new_n1093), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1100), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1097), .A2(new_n1099), .A3(KEYINPUT60), .A4(new_n602), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1107), .A2(new_n1092), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  INV_X1    g699(.A(G1996), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n995), .A2(new_n1125), .A3(new_n975), .A4(new_n983), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1129), .B2(new_n549), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n733), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1123), .A2(new_n1110), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1109), .B1(new_n1122), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1039), .B1(new_n1077), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1025), .B(new_n1135), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n999), .A2(new_n688), .B1(new_n684), .B2(new_n1091), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1008), .B1(new_n1137), .B2(new_n1016), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1001), .A2(G8), .A3(new_n1009), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1029), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1009), .B1(new_n1001), .B2(G8), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1010), .A2(new_n1143), .A3(new_n1038), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1144), .B2(new_n1026), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT127), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1132), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1123), .A2(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1108), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(new_n1057), .C1(new_n1052), .C2(new_n1063), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1149), .A2(new_n1151), .B1(KEYINPUT63), .B2(new_n1038), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1001), .A2(G8), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1008), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1037), .A3(new_n1139), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT63), .B1(new_n1157), .B2(new_n1025), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .A4(new_n1029), .ZN(new_n1160));
  OAI21_X1  g735(.A(G171), .B1(new_n1150), .B2(KEYINPUT62), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(KEYINPUT62), .B2(new_n1150), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1063), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1153), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1146), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT108), .ZN(new_n1166));
  OR3_X1    g741(.A1(new_n969), .A2(KEYINPUT107), .A3(new_n961), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT107), .B1(new_n969), .B2(new_n961), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1169), .A2(G1996), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n773), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(KEYINPUT108), .A3(new_n773), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n740), .B(new_n746), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1172), .B2(G1996), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1173), .B(new_n1174), .C1(new_n1169), .C2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT109), .Z(new_n1179));
  XNOR2_X1  g754(.A(new_n713), .B(new_n716), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1169), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1169), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(G1986), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1165), .A2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1169), .A2(G1986), .A3(G290), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT48), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1181), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n713), .A2(new_n715), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1179), .A2(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n740), .A2(G2067), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1169), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1170), .A2(KEYINPUT46), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1182), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1170), .A2(KEYINPUT46), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT47), .Z(new_n1197));
  NOR3_X1   g772(.A1(new_n1188), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G227), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n641), .B(new_n1201), .C1(new_n870), .C2(new_n872), .ZN(new_n1202));
  NOR3_X1   g776(.A1(new_n955), .A2(new_n956), .A3(new_n462), .ZN(new_n1203));
  INV_X1    g777(.A(G229), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1202), .A2(new_n1205), .ZN(G308));
  AOI21_X1  g780(.A(G401), .B1(new_n879), .B2(new_n882), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n1207), .A2(new_n1201), .A3(new_n1204), .A4(new_n1203), .ZN(G225));
endmodule


