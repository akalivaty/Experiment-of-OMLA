//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n450, new_n451, new_n453, new_n454,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G234));
  INV_X1    g027(.A(G2106), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G325));
  XOR2_X1   g035(.A(new_n459), .B(KEYINPUT68), .Z(G261));
  OAI22_X1  g036(.A1(new_n457), .A2(new_n453), .B1(new_n450), .B2(new_n458), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G101), .A3(G2104), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n467), .A2(new_n468), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(G136), .B2(new_n476), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT70), .Z(G162));
  OR2_X1    g062(.A1(new_n473), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n493), .A2(new_n494), .B1(G126), .B2(G2105), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n491), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n476), .B2(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT73), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(new_n502), .A3(KEYINPUT5), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n510), .B2(new_n511), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT75), .B(G51), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT72), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT72), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT6), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n516), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(KEYINPUT74), .A3(new_n528), .ZN(new_n529));
  AND4_X1   g104(.A1(G543), .A2(new_n523), .A3(new_n524), .A4(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n508), .A2(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n527), .A2(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT76), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n502), .B1(new_n536), .B2(new_n520), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(new_n524), .A3(new_n529), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n505), .A2(new_n507), .ZN(new_n544));
  INV_X1    g119(.A(new_n503), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n517), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G89), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n543), .A2(new_n548), .A3(new_n549), .A4(new_n535), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n541), .A2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n513), .B1(new_n537), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n542), .A2(G52), .A3(new_n529), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n513), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n542), .A2(G43), .A3(new_n529), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n547), .A2(G81), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT77), .Z(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND4_X1  g147(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n529), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n542), .A2(new_n575), .A3(G53), .A4(new_n529), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n547), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  NAND3_X1  g156(.A1(new_n557), .A2(KEYINPUT78), .A3(new_n558), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n542), .A2(G52), .A3(new_n529), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n556), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(G301));
  INV_X1    g161(.A(G166), .ZN(G303));
  NAND4_X1  g162(.A1(new_n523), .A2(G49), .A3(G543), .A4(new_n529), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n542), .A2(KEYINPUT79), .A3(G49), .A4(new_n529), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n537), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT80), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n592), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n598), .A2(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n513), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n508), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n517), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  AND3_X1   g182(.A1(new_n542), .A2(G47), .A3(new_n529), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n609), .A2(new_n513), .B1(new_n537), .B2(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n608), .A2(new_n611), .ZN(G290));
  AND2_X1   g187(.A1(new_n542), .A2(new_n529), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G54), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G651), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n537), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n614), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n582), .A2(new_n585), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G284));
  AOI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g204(.A(new_n628), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(new_n623), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n565), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n623), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n473), .A2(G2104), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n498), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  INV_X1    g220(.A(new_n481), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n646), .A2(G123), .B1(G135), .B2(new_n476), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n649));
  INV_X1    g224(.A(G111), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n649), .B2(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n644), .A2(new_n645), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT83), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n676), .B2(KEYINPUT18), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n654), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT84), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n688), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT85), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n689), .A2(new_n694), .A3(new_n691), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT86), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  NOR2_X1   g280(.A1(G29), .A2(G35), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G162), .B2(G29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT29), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2090), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n710), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n709), .B1(G1966), .B2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(G1966), .ZN(new_n714));
  NOR2_X1   g289(.A1(G171), .A2(new_n710), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G5), .B2(new_n710), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G1961), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G28), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OR2_X1    g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  NAND2_X1  g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  INV_X1    g300(.A(G129), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n481), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n476), .A2(G141), .ZN(new_n728));
  INV_X1    g303(.A(G105), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n639), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n720), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n720), .B2(G32), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n723), .B1(new_n720), .B2(new_n653), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n720), .B1(new_n736), .B2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G160), .B2(G29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n720), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n720), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n718), .A2(new_n735), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n720), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n646), .A2(G128), .B1(G140), .B2(new_n476), .ZN(new_n748));
  OR2_X1    g323(.A1(G104), .A2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT93), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G1961), .B2(new_n717), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n713), .A2(new_n714), .A3(new_n745), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n710), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n631), .B2(new_n710), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G19), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n566), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1341), .Z(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  INV_X1    g341(.A(new_n761), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n720), .A2(G33), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT94), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n476), .A2(G139), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n772), .B(new_n773), .C1(new_n473), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n733), .A2(new_n734), .B1(G2084), .B2(new_n739), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n762), .B(new_n768), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n710), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n577), .A2(new_n580), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n710), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n784), .B(new_n790), .C1(new_n783), .C2(new_n782), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n759), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(KEYINPUT89), .B1(new_n592), .B2(new_n596), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT89), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n795), .B(new_n595), .C1(new_n590), .C2(new_n591), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G16), .B2(G23), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT33), .B(G1976), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n799), .A2(new_n801), .ZN(new_n803));
  NOR2_X1   g378(.A1(G6), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n606), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  INV_X1    g381(.A(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n710), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n710), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT90), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1971), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n720), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n646), .A2(G119), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n476), .A2(G131), .ZN(new_n817));
  OR2_X1    g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n720), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  NAND2_X1  g399(.A1(G290), .A2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G24), .ZN(new_n826));
  OR3_X1    g401(.A1(new_n826), .A2(KEYINPUT87), .A3(G16), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT87), .B1(new_n826), .B2(G16), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT88), .B(G1986), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n814), .A2(new_n824), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT91), .B1(new_n813), .B2(KEYINPUT34), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n813), .A2(KEYINPUT91), .A3(KEYINPUT34), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n832), .B(new_n837), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n793), .B1(new_n836), .B2(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n792), .ZN(G150));
  NAND2_X1  g416(.A1(new_n613), .A2(G55), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n508), .A2(G67), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n513), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n845), .A2(KEYINPUT98), .B1(G93), .B2(new_n547), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n512), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n842), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(new_n565), .A3(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(new_n563), .ZN(new_n853));
  INV_X1    g428(.A(G81), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n561), .A2(new_n513), .B1(new_n537), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT99), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n613), .A2(G55), .B1(new_n848), .B2(new_n849), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n562), .A2(new_n563), .A3(new_n858), .A4(new_n564), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n846), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT38), .Z(new_n862));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n632), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n851), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  NAND2_X1  g445(.A1(new_n476), .A2(G142), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n875), .B2(G2105), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n646), .B2(G130), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n641), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n820), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G164), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n753), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n753), .A2(new_n883), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n885), .A2(new_n886), .B1(new_n730), .B2(new_n727), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n884), .A3(new_n731), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n889), .A3(new_n775), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n776), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n882), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n889), .ZN(new_n894));
  INV_X1    g469(.A(new_n776), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n881), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n880), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n898), .A3(new_n890), .ZN(new_n899));
  XNOR2_X1  g474(.A(G162), .B(G160), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n653), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n893), .A2(new_n899), .A3(KEYINPUT103), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n893), .B2(new_n899), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n851), .A2(new_n634), .ZN(new_n911));
  XNOR2_X1  g486(.A(G290), .B(G303), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n606), .B1(new_n794), .B2(new_n796), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n794), .A2(new_n796), .A3(new_n606), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n912), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(KEYINPUT105), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n861), .B(new_n636), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n631), .B1(KEYINPUT104), .B2(G299), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n787), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n631), .A2(new_n787), .A3(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n623), .B1(new_n787), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n928), .B2(new_n787), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n927), .A2(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n933), .B1(new_n926), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n925), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n911), .B1(new_n942), .B2(new_n634), .ZN(G295));
  OAI21_X1  g518(.A(new_n911), .B1(new_n942), .B2(new_n634), .ZN(G331));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n559), .A2(new_n540), .A3(new_n550), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n582), .A2(new_n585), .B1(new_n540), .B2(new_n550), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n861), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(new_n852), .A3(new_n860), .A4(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n935), .A2(new_n952), .A3(new_n939), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(new_n951), .A3(new_n937), .A4(new_n938), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n920), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n932), .A2(new_n960), .A3(new_n951), .A4(new_n949), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n953), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n921), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n955), .A2(new_n956), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n920), .B1(new_n953), .B2(new_n954), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n945), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n958), .B1(new_n957), .B2(new_n963), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(new_n945), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n967), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR4_X1   g552(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT108), .A4(new_n945), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n499), .B2(new_n500), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT109), .B(G40), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n472), .A2(new_n477), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n753), .B(G2067), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n731), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n988), .A2(G1996), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n991), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n731), .B(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n989), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n820), .B(new_n823), .Z(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n988), .ZN(new_n1002));
  OR2_X1    g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n987), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(KEYINPUT48), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(KEYINPUT48), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n821), .A2(new_n823), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n999), .A2(new_n1009), .B1(G2067), .B2(new_n754), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n987), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n997), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n797), .A2(G1976), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n1015));
  OAI21_X1  g590(.A(G125), .B1(new_n496), .B2(new_n497), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n473), .B1(new_n1016), .B2(new_n470), .ZN(new_n1017));
  OAI211_X1 g592(.A(G137), .B(new_n473), .C1(new_n496), .C2(new_n497), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n474), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1017), .A2(new_n1019), .A3(new_n984), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n473), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(G138), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G126), .A2(G2105), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1023), .A2(new_n480), .B1(new_n488), .B2(new_n490), .ZN(new_n1024));
  OAI211_X1 g599(.A(G138), .B(new_n473), .C1(new_n496), .C2(new_n497), .ZN(new_n1025));
  INV_X1    g600(.A(new_n494), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n598), .A2(new_n1032), .A3(new_n600), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1014), .A2(new_n1015), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n606), .A2(new_n807), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n603), .B2(new_n605), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT49), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1030), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n986), .B1(KEYINPUT45), .B2(new_n1028), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n981), .A2(KEYINPUT112), .A3(new_n982), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1971), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n986), .B1(new_n1048), .B2(new_n1028), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1028), .A2(KEYINPUT113), .A3(new_n1048), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(G2090), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n514), .B2(new_n518), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT55), .Z(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n794), .A2(new_n796), .A3(new_n1032), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT52), .B1(new_n1058), .B2(new_n1030), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1034), .A2(new_n1040), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1048), .B(new_n980), .C1(new_n499), .C2(new_n500), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1020), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1028), .A2(new_n1048), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1047), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT114), .B1(new_n1068), .B2(new_n1056), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1046), .A2(new_n1045), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(new_n1071), .C1(new_n1072), .C2(new_n1061), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2084), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1041), .A2(new_n983), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1061), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G168), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1060), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT115), .B1(new_n1082), .B2(KEYINPUT63), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1033), .A2(new_n1015), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1058), .A2(new_n1030), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1039), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1084), .B(new_n1085), .C1(new_n1090), .C2(new_n1081), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1056), .B1(G8), .B2(new_n1054), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(G168), .A3(KEYINPUT63), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1060), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1083), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1045), .B2(G2078), .ZN(new_n1097));
  INV_X1    g672(.A(G1961), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1053), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1096), .A2(G2078), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1097), .B(new_n1099), .C1(new_n1077), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n625), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1090), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n540), .A2(new_n550), .A3(KEYINPUT122), .A4(G8), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n540), .A2(new_n550), .A3(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT113), .B1(new_n1028), .B2(new_n1048), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n981), .A2(new_n1050), .A3(KEYINPUT50), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1063), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1112), .A2(new_n1075), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1106), .B(new_n1109), .C1(new_n1113), .C2(new_n1061), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1105), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1109), .A2(new_n1106), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1080), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1104), .A4(KEYINPUT51), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1109), .A2(new_n1106), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1120), .A2(KEYINPUT123), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT123), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(KEYINPUT62), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1119), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1103), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1032), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1035), .B1(new_n1130), .B2(G288), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1031), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1088), .A2(new_n1059), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1057), .ZN(new_n1134));
  INV_X1    g709(.A(G40), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n478), .A2(new_n1135), .A3(new_n1100), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n983), .A3(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1097), .A2(new_n1099), .A3(new_n1138), .ZN(new_n1139));
  OAI221_X1 g714(.A(KEYINPUT54), .B1(new_n1101), .B2(new_n625), .C1(new_n559), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1090), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1097), .A2(new_n1099), .A3(G301), .A4(new_n1138), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n625), .A2(new_n1101), .B1(new_n1143), .B2(KEYINPUT125), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1143), .A2(KEYINPUT125), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n789), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT117), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n536), .A2(G91), .A3(new_n508), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT116), .B(new_n1151), .C1(new_n578), .C2(new_n616), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n577), .A2(new_n1154), .A3(new_n580), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n577), .B2(new_n580), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1147), .B(new_n1150), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1147), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n577), .A2(new_n1154), .A3(new_n580), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1154), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G299), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1164));
  NOR2_X1   g739(.A1(new_n1029), .A2(G2067), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1053), .B2(new_n766), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n623), .B1(new_n1166), .B2(KEYINPUT60), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1165), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1112), .B2(G1348), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1163), .A2(new_n1164), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT118), .B(G1996), .Z(new_n1173));
  NAND4_X1  g748(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT58), .B(G1341), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1029), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1029), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1180), .A2(KEYINPUT59), .A3(new_n566), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT60), .B(new_n1168), .C1(new_n1112), .C2(G1348), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n631), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT59), .B1(new_n1180), .B2(new_n566), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT121), .B1(new_n1163), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1157), .A2(new_n1162), .A3(new_n1188), .A4(KEYINPUT61), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1172), .A2(new_n1185), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1162), .B1(new_n623), .B2(new_n1166), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1157), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1146), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1134), .B1(new_n1142), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1095), .A2(new_n1129), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(G290), .A2(G1986), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT111), .Z(new_n1197));
  INV_X1    g772(.A(new_n1004), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1001), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n987), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1195), .A2(KEYINPUT126), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT126), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1013), .B1(new_n1201), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g778(.A(G319), .ZN(new_n1205));
  OR3_X1    g779(.A1(G401), .A2(new_n1205), .A3(G227), .ZN(new_n1206));
  NOR2_X1   g780(.A1(G229), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g781(.A(new_n1207), .B(new_n909), .C1(new_n970), .C2(new_n966), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


