//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G43gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n210), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n208), .A2(G43gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n217), .A2(new_n218), .A3(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT14), .B(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n214), .B1(new_n213), .B2(new_n215), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n219), .B1(new_n229), .B2(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  INV_X1    g031(.A(G15gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(G22gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G15gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(G1gat), .B1(new_n234), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(G8gat), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n234), .A2(new_n236), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n237), .C1(new_n242), .C2(G1gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT89), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n228), .A2(new_n230), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n230), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT17), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n240), .A2(new_n243), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n253), .A3(new_n230), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT88), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n249), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n217), .A2(new_n218), .A3(new_n215), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n213), .A2(new_n215), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT87), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(new_n227), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n226), .B1(new_n216), .B2(new_n219), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n252), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT91), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n269), .A3(new_n252), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n257), .B(KEYINPUT13), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n271), .A2(KEYINPUT92), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT92), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n261), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n260), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT90), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n279), .A3(new_n260), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n206), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n206), .B1(new_n259), .B2(new_n260), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n261), .B(new_n283), .C1(new_n274), .C2(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT35), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT31), .B(G50gat), .ZN(new_n288));
  INV_X1    g087(.A(G106gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(G197gat), .ZN(new_n293));
  INV_X1    g092(.A(G204gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G197gat), .A2(G204gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(new_n297), .B2(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n308), .A2(KEYINPUT2), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n314), .A3(new_n308), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT76), .B(new_n312), .C1(new_n307), .C2(new_n309), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G228gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n303), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT3), .B1(new_n316), .B2(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT81), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n297), .A2(new_n299), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n302), .B1(new_n297), .B2(new_n299), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n305), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n323), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n320), .A2(new_n335), .A3(new_n323), .A4(new_n326), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G22gat), .ZN(new_n338));
  INV_X1    g137(.A(G78gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n328), .A2(new_n334), .A3(new_n235), .A4(new_n336), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n291), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G78gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n290), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT34), .ZN(new_n348));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT26), .ZN(new_n355));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n351), .A3(new_n350), .ZN(new_n363));
  AND4_X1   g162(.A1(new_n349), .A2(new_n353), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G183gat), .B2(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  OR3_X1    g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n370));
  NOR2_X1   g169(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n371));
  OAI22_X1  g170(.A1(new_n370), .A2(new_n371), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n358), .A2(new_n359), .B1(KEYINPUT23), .B2(new_n354), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n369), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n373), .B(KEYINPUT68), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(KEYINPUT25), .ZN(new_n379));
  INV_X1    g178(.A(new_n368), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n366), .B1(KEYINPUT69), .B2(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(KEYINPUT69), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n364), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G113gat), .B(G120gat), .Z(new_n386));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT72), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n396), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n389), .B(new_n390), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n402), .B2(new_n388), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n375), .A2(new_n376), .B1(new_n378), .B2(new_n383), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n364), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G227gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n322), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n348), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT34), .B(new_n409), .C1(new_n400), .C2(new_n406), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G15gat), .B(G43gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n406), .A3(new_n409), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n418), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n420), .B1(new_n411), .B2(new_n412), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n420), .A2(new_n411), .A3(new_n412), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n428), .A2(new_n429), .B1(new_n424), .B2(new_n423), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n343), .A2(new_n347), .A3(new_n427), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n287), .B1(new_n431), .B2(KEYINPUT85), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n343), .A2(new_n347), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n395), .A2(new_n318), .A3(new_n396), .A4(new_n398), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(KEYINPUT4), .B2(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n440));
  INV_X1    g239(.A(new_n325), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n399), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n435), .A2(new_n434), .A3(new_n437), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n439), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n319), .B1(new_n401), .B2(new_n403), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n443), .B1(new_n447), .B2(new_n435), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n446), .A2(new_n450), .A3(KEYINPUT5), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n404), .A2(new_n318), .A3(new_n437), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n442), .A2(new_n443), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT5), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n451), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT5), .B1(new_n448), .B2(new_n449), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n458), .B1(new_n471), .B2(new_n446), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n466), .B1(new_n472), .B2(new_n464), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n465), .B(new_n458), .C1(new_n471), .C2(new_n446), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n324), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n385), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT74), .B1(new_n405), .B2(new_n364), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n302), .ZN(new_n484));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT75), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n385), .B2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(new_n485), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT75), .B(new_n489), .C1(new_n405), .C2(new_n364), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n480), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n485), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n385), .A2(KEYINPUT29), .A3(new_n489), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n480), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n479), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n491), .B1(new_n485), .B2(new_n484), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n478), .C1(new_n499), .C2(new_n480), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n492), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n324), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n496), .A4(new_n478), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n425), .B1(new_n422), .B2(new_n426), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n433), .A2(new_n475), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n432), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n343), .A2(new_n347), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n501), .A2(new_n505), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n453), .A2(new_n455), .A3(new_n442), .ZN(new_n514));
  INV_X1    g313(.A(new_n443), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(new_n464), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n447), .A2(new_n435), .A3(new_n443), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT39), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n518), .B(new_n521), .C1(KEYINPUT83), .C2(KEYINPUT40), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n524), .B(new_n525), .C1(new_n464), .C2(new_n472), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n512), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n468), .B(new_n500), .C1(new_n473), .C2(new_n474), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n531), .B(new_n496), .C1(new_n499), .C2(new_n480), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n503), .A2(new_n534), .A3(new_n531), .A4(new_n496), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n478), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n494), .ZN(new_n537));
  INV_X1    g336(.A(new_n495), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n531), .B1(new_n539), .B2(new_n324), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n502), .A2(new_n480), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT38), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT37), .B1(new_n493), .B2(new_n497), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n536), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n528), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n475), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n512), .B1(new_n549), .B2(new_n513), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n507), .B2(new_n508), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n430), .A2(KEYINPUT36), .A3(new_n427), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n286), .B1(new_n511), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G190gat), .B(G218gat), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT7), .ZN(new_n564));
  OR2_X1    g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT97), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n566), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT97), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n574), .A2(new_n564), .A3(new_n567), .A4(new_n570), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n562), .B1(new_n250), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT98), .Z(new_n581));
  NAND3_X1  g380(.A1(new_n251), .A2(new_n254), .A3(new_n579), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n561), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n561), .A3(new_n582), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n559), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  INV_X1    g386(.A(new_n559), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G57gat), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n594), .A2(G64gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(G64gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G71gat), .B(G78gat), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n597), .ZN(new_n602));
  NOR2_X1   g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(KEYINPUT93), .B2(new_n591), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(KEYINPUT93), .B2(new_n591), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n244), .B1(new_n607), .B2(KEYINPUT21), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT95), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n609), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n600), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n602), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n602), .A2(new_n605), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n614), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n590), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n578), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n576), .B(new_n577), .C1(new_n601), .C2(new_n606), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n607), .A2(new_n578), .A3(KEYINPUT10), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n629), .ZN(new_n636));
  INV_X1    g435(.A(new_n630), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT100), .B(new_n628), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n628), .B1(new_n636), .B2(new_n637), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n632), .A2(new_n646), .A3(new_n633), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n632), .B2(new_n633), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n647), .A2(new_n648), .A3(new_n628), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n641), .A2(new_n638), .A3(new_n645), .ZN(new_n650));
  OAI22_X1  g449(.A1(new_n642), .A2(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n556), .A2(new_n626), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n475), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n231), .ZN(G1324gat));
  OR2_X1    g454(.A1(new_n653), .A2(new_n506), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(G8gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT42), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT42), .B2(new_n659), .ZN(G1325gat));
  NOR2_X1   g460(.A1(new_n554), .A2(KEYINPUT101), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n552), .B2(new_n553), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n653), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n509), .A2(new_n233), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n653), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n433), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n625), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n651), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n556), .A2(new_n590), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G29gat), .A3(new_n475), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT45), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n665), .A2(new_n548), .A3(new_n550), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n511), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n590), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  INV_X1    g480(.A(new_n590), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n511), .B2(new_n555), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  INV_X1    g484(.A(new_n206), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n259), .A2(new_n260), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n246), .A2(new_n248), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n268), .A2(new_n270), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n273), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT92), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n271), .A2(KEYINPUT92), .A3(new_n273), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n687), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n259), .A2(new_n279), .A3(new_n260), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n279), .B1(new_n259), .B2(new_n260), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n686), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n284), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n685), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n282), .A2(KEYINPUT102), .A3(new_n284), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n672), .A3(new_n651), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n684), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n221), .B1(new_n704), .B2(new_n549), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n676), .A2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n225), .B1(new_n707), .B2(KEYINPUT104), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n674), .A2(new_n506), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n704), .A2(new_n513), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G36gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n509), .A2(new_n211), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n674), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT106), .Z(new_n721));
  INV_X1    g520(.A(new_n665), .ZN(new_n722));
  INV_X1    g521(.A(new_n679), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n682), .B(new_n723), .C1(new_n677), .C2(new_n511), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n511), .A2(new_n555), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n681), .B1(new_n725), .B2(new_n590), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n722), .B(new_n703), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n718), .B1(new_n721), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n674), .B2(new_n719), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n211), .B1(new_n727), .B2(KEYINPUT107), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n684), .A2(new_n732), .A3(new_n722), .A4(new_n703), .ZN(new_n733));
  AOI211_X1 g532(.A(KEYINPUT108), .B(new_n730), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n733), .A3(G43gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n730), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n729), .B1(new_n734), .B2(new_n739), .ZN(G1330gat));
  NAND3_X1  g539(.A1(new_n684), .A2(new_n512), .A3(new_n703), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT48), .B1(new_n742), .B2(KEYINPUT109), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n674), .A2(G50gat), .A3(new_n433), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n742), .B(new_n744), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1331gat));
  INV_X1    g547(.A(new_n678), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n626), .A2(new_n702), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n652), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT110), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n678), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n475), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(new_n594), .ZN(G1332gat));
  OAI22_X1  g557(.A1(new_n756), .A2(new_n506), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT49), .B(G64gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n753), .A2(new_n513), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n753), .A2(new_n509), .A3(new_n755), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n768), .A3(new_n509), .A4(new_n755), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n753), .A2(G71gat), .A3(new_n722), .A4(new_n755), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT50), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1334gat));
  NOR2_X1   g575(.A1(new_n756), .A2(new_n433), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n339), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n702), .A2(new_n625), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT113), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n749), .A2(new_n682), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n549), .A2(new_n568), .A3(new_n651), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n780), .A2(new_n652), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n684), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n549), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n784), .A2(new_n785), .B1(new_n788), .B2(new_n568), .ZN(G1336gat));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n684), .A2(new_n513), .A3(new_n786), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n513), .A2(new_n569), .A3(new_n651), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n790), .B(new_n792), .C1(new_n784), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n782), .B2(new_n783), .ZN(new_n795));
  INV_X1    g594(.A(new_n792), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1337gat));
  NAND2_X1  g597(.A1(new_n787), .A2(new_n722), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G99gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n509), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n801), .A2(G99gat), .A3(new_n652), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n784), .B2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n684), .A2(new_n512), .A3(new_n786), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n512), .A2(new_n289), .A3(new_n651), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(new_n806), .C1(new_n784), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n782), .B2(new_n783), .ZN(new_n809));
  INV_X1    g608(.A(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n750), .A2(new_n651), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n632), .A2(new_n628), .A3(new_n633), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT54), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n632), .A2(new_n633), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n628), .B1(new_n818), .B2(KEYINPUT99), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n632), .A2(new_n646), .A3(new_n633), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n645), .B1(new_n634), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n815), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n649), .A2(new_n650), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT55), .B(new_n823), .C1(new_n649), .C2(new_n817), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n590), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n258), .B1(new_n249), .B2(new_n255), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n831), .A2(new_n832), .B1(new_n271), .B2(new_n273), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n205), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n284), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n700), .A2(new_n701), .A3(new_n829), .ZN(new_n838));
  INV_X1    g637(.A(new_n836), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n651), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n590), .B1(new_n841), .B2(KEYINPUT115), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n814), .B1(new_n845), .B2(new_n672), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n512), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(new_n549), .A3(new_n506), .A4(new_n509), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n286), .ZN(new_n850));
  NOR4_X1   g649(.A1(new_n847), .A2(new_n475), .A3(new_n513), .A4(new_n431), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n702), .A2(G113gat), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n849), .B2(new_n652), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n652), .A2(G120gat), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n849), .B2(new_n625), .ZN(new_n861));
  INV_X1    g660(.A(G127gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n862), .A3(new_n672), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1342gat));
  OAI21_X1  g663(.A(G134gat), .B1(new_n849), .B2(new_n682), .ZN(new_n865));
  INV_X1    g664(.A(new_n431), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n682), .A2(new_n513), .A3(G134gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n846), .A2(new_n549), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n722), .A2(new_n433), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n549), .A3(new_n872), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n873), .A2(G141gat), .A3(new_n513), .A4(new_n286), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n549), .A2(new_n506), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n722), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n846), .B2(new_n512), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n433), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n828), .B1(new_n282), .B2(new_n284), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n652), .A2(new_n836), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n285), .A2(new_n829), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n840), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n887), .A3(new_n682), .ZN(new_n888));
  INV_X1    g687(.A(new_n837), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n625), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n672), .B1(new_n888), .B2(new_n889), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n813), .B1(new_n894), .B2(KEYINPUT119), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n881), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n285), .B(new_n877), .C1(new_n878), .C2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n897), .A2(new_n898), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n875), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n702), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(new_n877), .C1(new_n878), .C2(new_n896), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n904), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT120), .B1(new_n904), .B2(G141gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(new_n874), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(G1344gat));
  INV_X1    g708(.A(new_n873), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n506), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n911), .A2(G148gat), .A3(new_n652), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n830), .A2(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n830), .A2(KEYINPUT123), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n839), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n888), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n625), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n626), .A2(new_n286), .A3(new_n652), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT57), .B(new_n433), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n879), .B1(new_n846), .B2(new_n512), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n877), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n652), .B1(new_n923), .B2(KEYINPUT122), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n922), .B(new_n924), .C1(KEYINPUT122), .C2(new_n923), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n913), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n913), .A2(G148gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n878), .A2(new_n896), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n923), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n929), .B2(new_n651), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n912), .B1(new_n926), .B2(new_n930), .ZN(G1345gat));
  NOR3_X1   g730(.A1(new_n911), .A2(KEYINPUT124), .A3(new_n625), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(G155gat), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n911), .B2(new_n625), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n672), .A2(G155gat), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT125), .Z(new_n936));
  AOI22_X1  g735(.A1(new_n933), .A2(new_n934), .B1(new_n929), .B2(new_n936), .ZN(G1346gat));
  INV_X1    g736(.A(G162gat), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n910), .A2(new_n938), .A3(new_n506), .A4(new_n590), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n928), .A2(new_n682), .A3(new_n923), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n938), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n847), .A2(new_n549), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n431), .A2(new_n506), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n903), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n848), .A2(new_n475), .A3(new_n513), .A4(new_n509), .ZN(new_n947));
  INV_X1    g746(.A(G169gat), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(new_n286), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n946), .A2(new_n949), .ZN(G1348gat));
  OAI21_X1  g749(.A(G176gat), .B1(new_n947), .B2(new_n652), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n652), .A2(G176gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n944), .B2(new_n952), .ZN(G1349gat));
  NAND3_X1  g752(.A1(new_n945), .A2(new_n350), .A3(new_n672), .ZN(new_n954));
  OAI21_X1  g753(.A(G183gat), .B1(new_n947), .B2(new_n625), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT60), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n351), .A3(new_n590), .ZN(new_n961));
  OAI21_X1  g760(.A(G190gat), .B1(new_n947), .B2(new_n682), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1351gat));
  NOR3_X1   g764(.A1(new_n722), .A2(new_n506), .A3(new_n433), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n942), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n293), .B1(new_n967), .B2(new_n702), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n722), .A2(new_n549), .A3(new_n506), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n922), .A2(G197gat), .A3(new_n285), .A4(new_n969), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(G1352gat));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n942), .A2(new_n294), .A3(new_n651), .A4(new_n966), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n922), .A2(new_n969), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n980), .B2(new_n652), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n979), .A3(new_n981), .ZN(G1353gat));
  OR3_X1    g781(.A1(new_n967), .A2(G211gat), .A3(new_n625), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n922), .A2(new_n672), .A3(new_n969), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n980), .A2(new_n988), .A3(new_n682), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n967), .B2(new_n682), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(G1355gat));
endmodule


