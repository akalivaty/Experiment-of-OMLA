//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955;
  XOR2_X1   g000(.A(KEYINPUT69), .B(G113gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT70), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n207), .C1(new_n204), .C2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G127gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G127gat), .B2(new_n210), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G127gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(KEYINPUT68), .C1(G127gat), .C2(new_n210), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n204), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n204), .A2(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n216), .B(new_n219), .C1(KEYINPUT68), .C2(new_n215), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT71), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT28), .Z(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n230), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n226), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  OAI21_X1  g036(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(new_n224), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n229), .B1(new_n233), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT65), .B(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n236), .B2(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n249), .B2(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n213), .A2(new_n220), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n222), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT64), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n252), .A2(new_n235), .A3(new_n253), .A4(new_n250), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT33), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G15gat), .B(G43gat), .Z(new_n263));
  XNOR2_X1  g062(.A(G71gat), .B(G99gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n259), .B(KEYINPUT32), .C1(new_n261), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n266), .B2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n258), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n256), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT34), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n257), .A2(KEYINPUT34), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n270), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT36), .ZN(new_n280));
  INV_X1    g079(.A(new_n278), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n281), .A2(new_n269), .A3(KEYINPUT72), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n272), .A2(new_n278), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(KEYINPUT72), .B2(new_n269), .ZN(new_n285));
  INV_X1    g084(.A(new_n282), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT36), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289));
  XNOR2_X1  g088(.A(G141gat), .B(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G155gat), .B(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n292), .B(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n290), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n297), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT79), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n304), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n305), .B(new_n252), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n252), .A2(new_n304), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT4), .ZN(new_n313));
  OR3_X1    g112(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n304), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n307), .B2(new_n221), .ZN(new_n318));
  INV_X1    g117(.A(new_n310), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT81), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n322), .A3(new_n314), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n311), .A3(new_n317), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(G57gat), .B(G85gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n321), .A2(new_n330), .A3(new_n325), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(KEYINPUT6), .A3(new_n331), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G226gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n251), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT73), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n346));
  OR2_X1    g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n345), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT74), .B1(new_n251), .B2(new_n340), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n251), .A2(KEYINPUT74), .A3(new_n340), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n343), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n251), .A2(new_n340), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n350), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  XOR2_X1   g155(.A(G8gat), .B(G36gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT75), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n354), .B2(new_n356), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n354), .A2(new_n368), .A3(new_n356), .A4(new_n361), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n289), .B1(new_n337), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n351), .B1(new_n305), .B2(new_n341), .ZN(new_n373));
  INV_X1    g172(.A(G228gat), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(new_n339), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n308), .B1(new_n350), .B2(KEYINPUT29), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n307), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n376), .A2(new_n304), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n379), .A2(new_n373), .B1(new_n374), .B2(new_n339), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G22gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT83), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT31), .B(G50gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n378), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(G22gat), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n383), .A2(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(KEYINPUT83), .A3(new_n389), .A4(new_n386), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n335), .A2(new_n336), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n366), .A2(new_n370), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT82), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n372), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n323), .A2(new_n309), .A3(new_n324), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n319), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT39), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n318), .A2(new_n319), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(KEYINPUT39), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n330), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT40), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(KEYINPUT40), .A3(new_n330), .A4(new_n404), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n332), .A4(new_n371), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n392), .A2(new_n394), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n354), .A2(new_n356), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n360), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT38), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n367), .A2(new_n369), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT38), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n353), .A2(new_n352), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n419), .A2(new_n351), .A3(new_n342), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n351), .B1(new_n355), .B2(new_n342), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n416), .B(new_n417), .C1(new_n423), .C2(new_n414), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n409), .B(new_n410), .C1(new_n424), .C2(new_n396), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n288), .A2(new_n399), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n410), .B1(new_n279), .B2(new_n282), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT35), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n396), .A2(new_n397), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n395), .B1(new_n285), .B2(new_n286), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n396), .A2(KEYINPUT82), .A3(new_n397), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT82), .B1(new_n396), .B2(new_n397), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n434), .B2(KEYINPUT35), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G78gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(G71gat), .A2(G78gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT9), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(G57gat), .A2(G64gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(G57gat), .A2(G64gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(G71gat), .A2(G78gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n438), .ZN(new_n447));
  AND2_X1   g246(.A1(G71gat), .A2(G78gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(G71gat), .A2(G78gat), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT94), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G57gat), .ZN(new_n453));
  INV_X1    g252(.A(G64gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(G57gat), .A3(G64gat), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n440), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n444), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT21), .ZN(new_n459));
  NAND2_X1  g258(.A1(G231gat), .A2(G233gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  XOR2_X1   g260(.A(G127gat), .B(G155gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT20), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n461), .B(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n465));
  XNOR2_X1  g264(.A(G183gat), .B(G211gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n464), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n382), .A2(G15gat), .ZN(new_n469));
  INV_X1    g268(.A(G15gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G22gat), .ZN(new_n471));
  INV_X1    g270(.A(G1gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT16), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(G1gat), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT89), .B1(new_n475), .B2(G1gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(G8gat), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  OAI221_X1 g278(.A(new_n474), .B1(KEYINPUT89), .B2(new_n479), .C1(G1gat), .C2(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n453), .A2(new_n454), .B1(new_n439), .B2(new_n438), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n447), .A3(new_n450), .A4(new_n456), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n443), .A2(new_n440), .ZN(new_n484));
  INV_X1    g283(.A(new_n437), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT96), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n489), .B2(KEYINPUT21), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n468), .B(new_n490), .Z(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n468), .B(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT41), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT99), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT100), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT105), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  INV_X1    g309(.A(G43gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(G50gat), .ZN(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G43gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n510), .B(KEYINPUT15), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n506), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n504), .A3(new_n505), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n504), .A2(new_n505), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n518), .A2(KEYINPUT86), .B1(new_n519), .B2(KEYINPUT14), .ZN(new_n520));
  NOR3_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT86), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT87), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NOR4_X1   g326(.A1(KEYINPUT86), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n516), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n518), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n506), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(new_n523), .A3(KEYINPUT87), .A4(new_n525), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n537), .B1(new_n546), .B2(new_n516), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n547), .B2(KEYINPUT17), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n540), .B(new_n537), .C1(new_n546), .C2(new_n516), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT101), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT101), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n552), .A2(new_n554), .A3(G85gat), .A4(G92gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT102), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G92gat), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT8), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT101), .B(new_n553), .C1(new_n560), .C2(new_n556), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n555), .A2(new_n561), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n562), .ZN(new_n566));
  NOR2_X1   g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT103), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT103), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n562), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n565), .A2(new_n572), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n550), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT104), .B1(new_n549), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n549), .A2(KEYINPUT104), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n499), .A2(KEYINPUT41), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n575), .B2(new_n547), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n503), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  AOI211_X1 g384(.A(KEYINPUT105), .B(new_n583), .C1(new_n579), .C2(new_n580), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n502), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n580), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT105), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n581), .A2(new_n503), .A3(new_n584), .ZN(new_n594));
  INV_X1    g393(.A(new_n502), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n587), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n590), .B1(new_n587), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n487), .B1(new_n573), .B2(new_n574), .ZN(new_n601));
  AND2_X1   g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n568), .A2(new_n571), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n555), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n565), .A2(new_n572), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n458), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n489), .A2(KEYINPUT10), .A3(new_n576), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n601), .A2(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT106), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT106), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n614), .B(KEYINPUT10), .C1(new_n601), .C2(new_n607), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n610), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n602), .B(KEYINPUT107), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n609), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  OR2_X1    g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n488), .A2(new_n612), .A3(new_n575), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n573), .A2(new_n574), .A3(new_n487), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n458), .B1(new_n605), .B2(new_n606), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n612), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n614), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n611), .A2(KEYINPUT106), .A3(new_n612), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n608), .B(new_n622), .C1(new_n630), .C2(new_n602), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n497), .A2(new_n600), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G197gat), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT11), .B(G169gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n539), .B(new_n481), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n547), .B1(new_n480), .B2(new_n478), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT90), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n481), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT90), .B1(new_n478), .B2(new_n480), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n550), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n646), .B1(new_n549), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n651), .B2(new_n642), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT18), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n642), .ZN(new_n655));
  AOI211_X1 g454(.A(new_n655), .B(new_n646), .C1(new_n549), .C2(new_n650), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(new_n645), .A3(KEYINPUT18), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n639), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT18), .B1(new_n656), .B2(new_n645), .ZN(new_n660));
  INV_X1    g459(.A(new_n639), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n644), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n634), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n436), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n337), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n371), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n671), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n479), .B1(new_n666), .B2(new_n371), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n673), .A2(new_n674), .B1(new_n669), .B2(new_n670), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT108), .B1(new_n671), .B2(KEYINPUT42), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n285), .A2(new_n286), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n666), .A2(new_n470), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n436), .A2(new_n288), .A3(new_n665), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n470), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n395), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  OAI21_X1  g483(.A(new_n599), .B1(new_n426), .B2(new_n435), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n497), .A2(new_n664), .A3(new_n632), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n504), .A3(new_n337), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n288), .A2(new_n399), .A3(new_n425), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n430), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n599), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n337), .A3(new_n687), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n698), .A2(KEYINPUT109), .A3(new_n337), .A4(new_n687), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(G29gat), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n691), .A2(new_n703), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n688), .A2(G36gat), .A3(new_n397), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT46), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n698), .A2(new_n371), .A3(new_n687), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n505), .B2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n288), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n697), .A3(new_n709), .A4(new_n687), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n511), .B1(new_n710), .B2(KEYINPUT110), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT110), .B2(new_n710), .ZN(new_n712));
  INV_X1    g511(.A(new_n678), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n688), .A2(G43gat), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n710), .A2(G43gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n718), .B2(new_n714), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n689), .A2(new_n513), .A3(new_n395), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n693), .A2(new_n697), .A3(new_n395), .A4(new_n687), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G50gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1331gat));
  NAND4_X1  g525(.A1(new_n497), .A2(new_n664), .A3(new_n600), .A4(new_n632), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n436), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n337), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n371), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n709), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n713), .A2(G71gat), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n735), .A2(G71gat), .B1(new_n728), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n728), .A2(new_n395), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n497), .A2(new_n663), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n599), .A4(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n599), .B(new_n741), .C1(new_n426), .C2(new_n435), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n749), .A2(new_n560), .A3(new_n337), .A4(new_n632), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n497), .A2(new_n663), .A3(new_n633), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n698), .A2(new_n337), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n560), .B2(new_n752), .ZN(G1336gat));
  NOR3_X1   g552(.A1(new_n397), .A2(G92gat), .A3(new_n633), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n693), .A2(new_n697), .A3(new_n371), .A4(new_n751), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n557), .A2(new_n559), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n748), .A2(new_n742), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n756), .A2(new_n757), .B1(new_n762), .B2(new_n754), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n755), .A2(new_n760), .B1(new_n761), .B2(new_n763), .ZN(G1337gat));
  INV_X1    g563(.A(G99gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n765), .A3(new_n678), .A4(new_n632), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n698), .A2(new_n709), .A3(new_n751), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1338gat));
  NOR3_X1   g567(.A1(new_n410), .A2(G106gat), .A3(new_n633), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT113), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n749), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n693), .A2(new_n697), .A3(new_n395), .A4(new_n751), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT53), .B1(new_n773), .B2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n773), .A2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n762), .B2(new_n771), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT114), .B(new_n770), .C1(new_n748), .C2(new_n742), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  NOR2_X1   g581(.A1(new_n634), .A2(new_n663), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n497), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n617), .B(new_n610), .C1(new_n613), .C2(new_n615), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT54), .B(new_n786), .C1(new_n630), .C2(new_n602), .ZN(new_n787));
  INV_X1    g586(.A(new_n622), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n616), .A2(new_n789), .A3(new_n618), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n631), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(KEYINPUT115), .A3(new_n631), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n651), .A2(new_n642), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n640), .A2(new_n643), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n638), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n662), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n799), .A2(new_n597), .A3(new_n598), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n794), .A2(new_n663), .A3(new_n795), .A4(new_n798), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n632), .A2(new_n662), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n599), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(KEYINPUT116), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n785), .B1(new_n811), .B2(KEYINPUT117), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813));
  AOI211_X1 g612(.A(new_n813), .B(new_n804), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n784), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n337), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n427), .A2(new_n371), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n663), .A2(new_n202), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n815), .A2(new_n410), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n713), .A2(new_n396), .A3(new_n371), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n664), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1340gat));
  NOR2_X1   g626(.A1(new_n633), .A2(G120gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n820), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G120gat), .B1(new_n825), .B2(new_n633), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n825), .B2(new_n785), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n785), .A2(G127gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n818), .B2(new_n833), .ZN(G1342gat));
  NAND3_X1  g633(.A1(new_n823), .A2(new_n599), .A3(new_n824), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G134gat), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n599), .A2(new_n214), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n817), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n816), .A2(new_n840), .A3(new_n817), .A4(new_n837), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n836), .A2(new_n839), .A3(KEYINPUT119), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(new_n287), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n285), .A2(KEYINPUT36), .A3(new_n286), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n395), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(new_n371), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n664), .A2(G141gat), .ZN(new_n853));
  AND4_X1   g652(.A1(new_n337), .A2(new_n852), .A3(new_n815), .A4(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n815), .A2(new_n855), .A3(new_n395), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n288), .A2(new_n337), .A3(new_n397), .ZN(new_n857));
  INV_X1    g656(.A(new_n804), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n798), .A2(new_n631), .A3(new_n791), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n806), .B1(new_n664), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n806), .B(KEYINPUT120), .C1(new_n664), .C2(new_n859), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n600), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n497), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n395), .B1(new_n865), .B2(new_n783), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n857), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n856), .A2(new_n663), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n854), .B1(new_n868), .B2(G141gat), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n868), .B2(G141gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  AOI221_X4 g672(.A(new_n854), .B1(new_n870), .B2(new_n873), .C1(G141gat), .C2(new_n868), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1344gat));
  AND2_X1   g674(.A1(new_n816), .A2(new_n852), .ZN(new_n876));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n632), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n856), .A2(new_n867), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n877), .C1(new_n879), .C2(new_n632), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n815), .A2(KEYINPUT57), .A3(new_n395), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n855), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n857), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n632), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n881), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n878), .B1(new_n880), .B2(new_n887), .ZN(G1345gat));
  NAND3_X1  g687(.A1(new_n876), .A2(new_n294), .A3(new_n497), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n879), .A2(new_n497), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n294), .ZN(G1346gat));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n295), .A3(new_n599), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n879), .A2(new_n599), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n295), .ZN(G1347gat));
  AND2_X1   g693(.A1(new_n815), .A2(new_n396), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n427), .A2(new_n397), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n895), .A2(new_n227), .A3(new_n663), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT123), .Z(new_n898));
  NAND2_X1  g697(.A1(new_n396), .A2(new_n371), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n713), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n823), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n664), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(G1348gat));
  INV_X1    g702(.A(new_n246), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n901), .A2(new_n904), .A3(new_n633), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n228), .B1(new_n906), .B2(new_n633), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT124), .B(new_n228), .C1(new_n906), .C2(new_n633), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1349gat));
  OAI21_X1  g710(.A(G183gat), .B1(new_n901), .B2(new_n785), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n223), .A3(new_n497), .A4(new_n896), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n901), .B2(new_n600), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n599), .A2(new_n224), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n920), .A2(new_n921), .B1(new_n906), .B2(new_n922), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n849), .A2(new_n397), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n895), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT125), .B(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n663), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n709), .A2(new_n899), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n882), .B2(new_n883), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(KEYINPUT126), .A3(new_n663), .ZN(new_n931));
  INV_X1    g730(.A(new_n926), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT126), .B1(new_n930), .B2(new_n663), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n633), .A2(G204gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n895), .A2(new_n924), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  INV_X1    g737(.A(new_n930), .ZN(new_n939));
  OAI21_X1  g738(.A(G204gat), .B1(new_n939), .B2(new_n633), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n937), .B2(KEYINPUT62), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n938), .B(new_n940), .C1(new_n942), .C2(new_n944), .ZN(G1353gat));
  INV_X1    g744(.A(G211gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n946), .A3(new_n497), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n497), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  AOI211_X1 g749(.A(new_n950), .B(new_n946), .C1(new_n930), .C2(new_n497), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n949), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n939), .B2(new_n600), .ZN(new_n953));
  INV_X1    g752(.A(G218gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n925), .A2(new_n954), .A3(new_n599), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1355gat));
endmodule


