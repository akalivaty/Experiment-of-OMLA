//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G50), .C2(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n203), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n206), .A2(G50), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT66), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(KEYINPUT66), .A3(G13), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n227), .B1(new_n221), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT8), .B(G58), .Z(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n262), .B1(new_n256), .B2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G58), .A2(G68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n204), .A2(new_n205), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G159), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(G20), .A3(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT72), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT72), .ZN(new_n272));
  AOI211_X1 g0072(.A(new_n272), .B(new_n269), .C1(new_n266), .C2(G20), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n257), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n253), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n253), .A4(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G68), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT16), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n203), .B1(new_n280), .B2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT16), .ZN(new_n286));
  NOR4_X1   g0086(.A1(new_n271), .A2(new_n273), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n264), .B1(new_n288), .B2(new_n258), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(G1), .B(G13), .C1(new_n257), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n290), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n218), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n276), .A2(new_n277), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G223), .B2(G1698), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G226), .ZN(new_n300));
  INV_X1    g0100(.A(G87), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n298), .A2(new_n300), .B1(new_n257), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n294), .ZN(new_n303));
  AOI211_X1 g0103(.A(new_n292), .B(new_n296), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(KEYINPUT74), .A2(G190), .ZN(new_n307));
  NAND2_X1  g0107(.A1(KEYINPUT74), .A2(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n289), .A2(KEYINPUT17), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n267), .A2(new_n270), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n272), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n270), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n283), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n286), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n274), .A2(KEYINPUT16), .A3(new_n283), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n258), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(new_n306), .A3(new_n263), .A4(new_n309), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n263), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n302), .A2(new_n303), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  INV_X1    g0124(.A(new_n292), .ZN(new_n325));
  INV_X1    g0125(.A(new_n296), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n304), .B2(G169), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n322), .A2(KEYINPUT18), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT18), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n289), .B2(new_n328), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n328), .B1(new_n317), .B2(new_n263), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n336), .A2(KEYINPUT73), .A3(KEYINPUT18), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n321), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n299), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n297), .B(new_n341), .C1(G232), .C2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n294), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n295), .A2(new_n219), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n292), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR4_X1   g0148(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT13), .A4(new_n292), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(G179), .B1(KEYINPUT71), .B2(KEYINPUT14), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT71), .B1(new_n352), .B2(KEYINPUT14), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G169), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(G169), .B(new_n353), .C1(new_n348), .C2(new_n349), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n257), .A2(G20), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n360));
  INV_X1    g0160(.A(G50), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G20), .A2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n258), .ZN(new_n365));
  XOR2_X1   g0165(.A(new_n365), .B(KEYINPUT11), .Z(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT68), .B1(new_n252), .B2(new_n255), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n252), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n369));
  INV_X1    g0169(.A(new_n258), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n368), .A2(new_n250), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n203), .B1(new_n371), .B2(KEYINPUT12), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n373), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n256), .A2(KEYINPUT12), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n366), .A2(new_n372), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n350), .A2(G190), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n376), .B(new_n379), .C1(new_n305), .C2(new_n350), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n339), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n259), .A2(G50), .A3(new_n250), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n252), .A2(new_n255), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n260), .A2(new_n359), .B1(G150), .B2(new_n362), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n382), .B1(G50), .B2(new_n383), .C1(new_n370), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  MUX2_X1   g0189(.A(G222), .B(G223), .S(G1698), .Z(new_n390));
  AND2_X1   g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(KEYINPUT3), .A2(G33), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n303), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n297), .A2(G77), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n325), .B1(new_n340), .B2(new_n295), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n387), .A2(new_n388), .B1(G200), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(KEYINPUT69), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n389), .A2(new_n397), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT10), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n355), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n396), .A2(G179), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n387), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(G232), .B(new_n299), .C1(new_n391), .C2(new_n392), .ZN(new_n408));
  OAI211_X1 g0208(.A(G238), .B(G1698), .C1(new_n391), .C2(new_n392), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n209), .C2(new_n297), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n292), .B1(new_n410), .B2(new_n303), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT67), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n294), .A2(G244), .A3(new_n290), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g0216(.A(G190), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n359), .ZN(new_n420));
  INV_X1    g0220(.A(G77), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n253), .B2(new_n421), .C1(new_n363), .C2(new_n261), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n258), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n373), .A2(new_n421), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(new_n421), .C2(new_n371), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n416), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G200), .A3(new_n414), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n417), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n414), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n324), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n355), .A3(new_n414), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n425), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n381), .A2(new_n407), .A3(new_n430), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  XOR2_X1   g0237(.A(G97), .B(G107), .Z(new_n438));
  INV_X1    g0238(.A(KEYINPUT6), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT75), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n439), .B2(new_n209), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(G97), .B(G107), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n440), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n445), .B1(new_n442), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g0247(.A(G20), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n282), .A2(G107), .B1(G77), .B2(new_n362), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n258), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n256), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n249), .A2(G33), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n259), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n297), .A2(G244), .A3(new_n299), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT77), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n460), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n297), .A2(G244), .A3(new_n299), .A4(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n303), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n291), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n294), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G257), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n467), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n355), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n466), .A2(new_n303), .B1(G257), .B2(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n324), .A3(new_n475), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n457), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n455), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n383), .A2(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT25), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT23), .B1(new_n253), .B2(G107), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT23), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n209), .A3(G20), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n253), .A2(G33), .A3(G116), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n253), .B(G87), .C1(new_n391), .C2(new_n392), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n297), .A2(KEYINPUT22), .A3(new_n253), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n488), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(new_n496), .ZN(new_n504));
  INV_X1    g0304(.A(new_n488), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n500), .A4(new_n501), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n487), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n484), .B(new_n486), .C1(new_n507), .C2(new_n370), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n477), .A2(KEYINPUT84), .A3(G264), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n476), .B2(new_n210), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n297), .A2(G257), .A3(G1698), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n297), .A2(G250), .A3(new_n299), .ZN(new_n513));
  INV_X1    g0313(.A(G294), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n257), .C2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n509), .A2(new_n511), .B1(new_n515), .B2(new_n303), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n475), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n355), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n324), .A3(new_n475), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n508), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n450), .A2(new_n258), .B1(new_n452), .B2(new_n256), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n479), .A2(G200), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n481), .A2(G190), .A3(new_n475), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n456), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n359), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n253), .B1(new_n343), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n301), .A2(new_n452), .A3(new_n209), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n297), .A2(new_n253), .A3(G68), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n258), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n383), .A2(G87), .A3(new_n370), .A4(new_n454), .ZN(new_n533));
  INV_X1    g0333(.A(new_n369), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n367), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n532), .B(new_n533), .C1(new_n535), .C2(new_n419), .ZN(new_n536));
  INV_X1    g0336(.A(G244), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G1698), .ZN(new_n538));
  OAI221_X1 g0338(.A(new_n538), .B1(G238), .B2(G1698), .C1(new_n391), .C2(new_n392), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n294), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n469), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n294), .A2(new_n542), .A3(G250), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n542), .A2(new_n291), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n305), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR4_X1   g0348(.A1(new_n541), .A2(new_n544), .A3(new_n398), .A4(new_n546), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n536), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n541), .A2(new_n546), .A3(new_n544), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT78), .B1(new_n551), .B2(new_n324), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n539), .A2(new_n540), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n303), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n324), .A3(new_n547), .A4(new_n543), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n551), .B2(G169), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n556), .B2(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n455), .A2(new_n419), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n373), .A2(new_n418), .B1(new_n258), .B2(new_n531), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n483), .A2(new_n520), .A3(new_n524), .A4(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(new_n299), .C1(new_n391), .C2(new_n392), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(G1698), .C1(new_n391), .C2(new_n392), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT79), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n303), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n474), .B1(new_n477), .B2(G270), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(KEYINPUT80), .A3(new_n303), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n535), .A2(G116), .A3(new_n370), .A4(new_n454), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n373), .A2(new_n214), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n462), .B(new_n253), .C1(G33), .C2(new_n452), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n258), .C1(new_n253), .C2(G116), .ZN(new_n580));
  XOR2_X1   g0380(.A(new_n580), .B(KEYINPUT20), .Z(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n576), .A2(G169), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n576), .A2(new_n585), .A3(G169), .A4(new_n582), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n573), .A2(G179), .A3(new_n574), .A4(new_n575), .ZN(new_n588));
  INV_X1    g0388(.A(new_n582), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT80), .B1(new_n570), .B2(new_n303), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n572), .B(new_n294), .C1(new_n567), .C2(new_n569), .ZN(new_n592));
  INV_X1    g0392(.A(new_n574), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(KEYINPUT81), .A3(G179), .A4(new_n582), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n584), .A2(new_n586), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n576), .A2(G200), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n307), .A2(new_n308), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n589), .C1(new_n598), .C2(new_n576), .ZN(new_n599));
  INV_X1    g0399(.A(new_n508), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n516), .A2(G190), .A3(new_n475), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n517), .A2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n562), .A2(new_n596), .A3(new_n599), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n437), .A2(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n406), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n334), .A2(new_n330), .ZN(new_n607));
  INV_X1    g0407(.A(new_n378), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n380), .B1(new_n608), .B2(new_n435), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n321), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n606), .B1(new_n610), .B2(new_n403), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n584), .A2(new_n586), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n590), .A2(new_n595), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n520), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT85), .B1(new_n536), .B2(new_n548), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n554), .A2(new_n547), .A3(new_n543), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n559), .A2(new_n617), .A3(new_n618), .A4(new_n533), .ZN(new_n619));
  INV_X1    g0419(.A(new_n549), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n603), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n483), .A2(new_n524), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n560), .B(new_n555), .C1(G169), .C2(new_n551), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(new_n483), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n561), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n621), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n483), .A3(KEYINPUT26), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n611), .B1(new_n437), .B2(new_n633), .ZN(G369));
  NOR2_X1   g0434(.A1(new_n251), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n249), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n520), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n612), .A2(new_n613), .A3(new_n599), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n582), .A2(new_n641), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n596), .B2(new_n644), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n596), .A2(new_n641), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n641), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n603), .B1(new_n600), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n520), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n642), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n642), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT86), .Z(G399));
  INV_X1    g0456(.A(new_n224), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n528), .A2(G116), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G1), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n230), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n627), .A2(new_n626), .A3(new_n561), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n629), .B2(new_n483), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n624), .A2(new_n666), .A3(new_n625), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n650), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(KEYINPUT29), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n632), .A2(new_n650), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(KEYINPUT29), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT30), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n591), .A2(new_n592), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n675), .A2(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(G179), .A3(new_n574), .A4(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n481), .A2(new_n475), .A3(new_n516), .A4(new_n551), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n591), .A2(new_n592), .A3(new_n324), .A4(new_n593), .ZN(new_n682));
  INV_X1    g0482(.A(new_n680), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n675), .A4(KEYINPUT30), .ZN(new_n684));
  AOI21_X1  g0484(.A(G179), .B1(new_n481), .B2(new_n475), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n576), .A2(new_n685), .A3(new_n517), .A4(new_n616), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT31), .B1(new_n687), .B2(new_n641), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n643), .A2(new_n603), .A3(new_n562), .A4(new_n650), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n673), .B(new_n674), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n641), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n604), .C2(new_n641), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT88), .B1(new_n697), .B2(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n672), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n663), .B1(new_n701), .B2(G1), .ZN(G364));
  NOR2_X1   g0502(.A1(G13), .A2(G33), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G20), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n646), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n251), .A2(new_n468), .A3(G20), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT89), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(new_n658), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT90), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n297), .A2(G355), .A3(new_n224), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n657), .A2(new_n297), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n246), .B2(new_n468), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n230), .A2(G45), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n715), .B1(G116), .B2(new_n224), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n227), .B1(G20), .B2(new_n355), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n705), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n253), .A2(G190), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n324), .A3(new_n305), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n268), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(KEYINPUT32), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n253), .A2(new_n324), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G200), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G190), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(G68), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n598), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G50), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n305), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n723), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n297), .B1(new_n736), .B2(new_n209), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n728), .A2(new_n305), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n598), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(G20), .A3(G190), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n202), .B1(new_n301), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n398), .A2(G179), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n253), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n737), .B(new_n742), .C1(G97), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n738), .A2(G190), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n726), .A2(KEYINPUT32), .B1(G77), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n732), .A2(new_n734), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n733), .A2(G326), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT33), .B(G317), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n750), .B1(new_n731), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n740), .A2(new_n753), .B1(new_n754), .B2(new_n741), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(G311), .B2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n736), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n297), .B1(new_n757), .B2(G283), .ZN(new_n758));
  INV_X1    g0558(.A(new_n724), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G329), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n752), .A2(new_n756), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n744), .A2(new_n514), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n749), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n720), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n707), .A2(new_n714), .A3(new_n722), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n647), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n712), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n646), .A2(G330), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT94), .Z(G396));
  NOR2_X1   g0571(.A1(new_n434), .A2(new_n641), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n425), .A2(new_n641), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n429), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n434), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n773), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n426), .B1(new_n324), .B2(new_n431), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(new_n433), .B1(new_n429), .B2(new_n775), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT96), .B1(new_n780), .B2(new_n772), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n670), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n699), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n632), .A2(new_n650), .A3(new_n782), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n785), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n712), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n757), .A2(G87), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n740), .B2(new_n514), .ZN(new_n792));
  INV_X1    g0592(.A(new_n741), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n297), .B(new_n792), .C1(G107), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n731), .A2(G283), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n745), .A2(G97), .B1(new_n759), .B2(G311), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n733), .A2(G303), .B1(G116), .B2(new_n747), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n731), .A2(G150), .B1(new_n733), .B2(G137), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  INV_X1    g0600(.A(new_n747), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n740), .C1(new_n268), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT34), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n741), .A2(new_n361), .B1(new_n736), .B2(new_n203), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G132), .B2(new_n759), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(new_n297), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n744), .A2(new_n202), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n720), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n720), .A2(new_n703), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n713), .B1(new_n421), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT95), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n809), .B(new_n812), .C1(new_n704), .C2(new_n782), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n790), .A2(new_n813), .ZN(G384));
  INV_X1    g0614(.A(KEYINPUT40), .ZN(new_n815));
  INV_X1    g0615(.A(new_n318), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n317), .A2(new_n263), .B1(new_n328), .B2(new_n639), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n816), .A2(KEYINPUT37), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  INV_X1    g0620(.A(new_n817), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n318), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT100), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT101), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT101), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT37), .B1(new_n816), .B2(new_n817), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(KEYINPUT100), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n819), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n639), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n322), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n607), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n321), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT101), .B1(new_n822), .B2(new_n823), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n826), .A2(KEYINPUT100), .A3(new_n825), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n818), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n828), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n339), .B2(new_n830), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n318), .B(KEYINPUT17), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT73), .B1(new_n336), .B2(KEYINPUT18), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n336), .A2(KEYINPUT18), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n337), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT99), .A3(new_n831), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n819), .A2(new_n826), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n841), .A2(new_n847), .A3(KEYINPUT38), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n839), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n377), .A2(new_n641), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n378), .A2(new_n380), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n358), .A2(new_n377), .A3(new_n641), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n782), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(new_n697), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n815), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n841), .A2(new_n848), .A3(new_n847), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n838), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n849), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n855), .A2(new_n697), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT102), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n674), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n695), .A2(new_n696), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n612), .A2(new_n613), .A3(new_n599), .A4(new_n603), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n520), .A2(new_n483), .A3(new_n561), .A4(new_n524), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(new_n641), .ZN(new_n871));
  OAI21_X1  g0671(.A(G330), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n437), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT103), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n697), .B1(new_n876), .B2(new_n857), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n437), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n378), .A2(new_n641), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n839), .A2(new_n882), .A3(new_n849), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n862), .A2(new_n849), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n786), .A2(new_n773), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n854), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n885), .A2(new_n887), .B1(new_n607), .B2(new_n829), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n878), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n436), .B1(new_n669), .B2(new_n671), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n611), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n249), .B2(new_n635), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n446), .A2(new_n447), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT98), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n214), .B1(new_n896), .B2(KEYINPUT35), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n227), .A2(new_n253), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(KEYINPUT35), .C2(new_n896), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n265), .A2(G77), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n230), .A2(new_n901), .B1(G50), .B2(new_n203), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n251), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(new_n900), .A3(new_n903), .ZN(G367));
  NAND4_X1  g0704(.A1(new_n653), .A2(new_n623), .A3(new_n614), .A4(new_n648), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT42), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n457), .A2(new_n641), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n623), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n483), .B1(new_n908), .B2(new_n520), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n650), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n536), .A2(new_n641), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n625), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n625), .A2(new_n621), .A3(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n906), .A2(new_n910), .B1(KEYINPUT43), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n767), .A2(new_n654), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n483), .B2(new_n650), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n917), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n658), .B(new_n922), .Z(new_n923));
  NOR2_X1   g0723(.A1(new_n520), .A2(new_n641), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n652), .B2(new_n648), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n919), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT44), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n919), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT45), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n918), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n649), .B(new_n653), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n701), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n931), .B1(new_n930), .B2(KEYINPUT105), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n923), .B1(new_n936), .B2(new_n701), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n711), .B(KEYINPUT106), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n921), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n914), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n713), .B1(new_n941), .B2(new_n705), .ZN(new_n942));
  INV_X1    g0742(.A(new_n716), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n721), .B1(new_n224), .B2(new_n418), .C1(new_n239), .C2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n731), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n945), .A2(new_n268), .B1(new_n361), .B2(new_n801), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(G137), .B2(new_n759), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n745), .A2(G68), .ZN(new_n949));
  INV_X1    g0749(.A(new_n733), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n949), .C1(new_n800), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n736), .A2(new_n421), .ZN(new_n952));
  INV_X1    g0752(.A(G150), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n740), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n946), .A2(new_n947), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n951), .A2(new_n952), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n297), .C1(new_n202), .C2(new_n741), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT108), .Z(new_n958));
  OAI21_X1  g0758(.A(new_n393), .B1(new_n736), .B2(new_n452), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT46), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n741), .B2(new_n214), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n724), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n959), .B(new_n963), .C1(G303), .C2(new_n739), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n733), .A2(G311), .B1(G283), .B2(new_n747), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n731), .A2(G294), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n741), .A2(new_n960), .A3(new_n214), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G107), .B2(new_n745), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n958), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  INV_X1    g0771(.A(new_n720), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n942), .B(new_n944), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n940), .A2(new_n973), .ZN(G387));
  NOR2_X1   g0774(.A1(new_n933), .A2(new_n701), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n934), .A2(new_n975), .A3(new_n659), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n933), .A2(new_n939), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT109), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n716), .B1(new_n236), .B2(new_n468), .ZN(new_n979));
  INV_X1    g0779(.A(new_n660), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n224), .A3(new_n297), .ZN(new_n981));
  AOI211_X1 g0781(.A(G45), .B(new_n980), .C1(G68), .C2(G77), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n260), .A2(new_n361), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT50), .Z(new_n984));
  AOI22_X1  g0784(.A1(new_n979), .A2(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n224), .A2(G107), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n721), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n714), .B(new_n987), .C1(new_n653), .C2(new_n706), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n731), .A2(G311), .B1(new_n733), .B2(G322), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n754), .B2(new_n801), .C1(new_n962), .C2(new_n740), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  INV_X1    g0791(.A(G283), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n992), .B2(new_n744), .C1(new_n514), .C2(new_n741), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT49), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G326), .A2(new_n759), .B1(new_n757), .B2(G116), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n393), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n744), .A2(new_n418), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n793), .A2(G77), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n953), .B2(new_n724), .C1(new_n950), .C2(new_n268), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G50), .C2(new_n739), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n203), .B2(new_n801), .C1(new_n261), .C2(new_n945), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n297), .B1(new_n736), .B2(new_n452), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n988), .B1(new_n1003), .B2(new_n720), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n976), .A2(new_n978), .A3(new_n1005), .ZN(G393));
  XNOR2_X1  g0806(.A(new_n930), .B(new_n918), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n936), .B(new_n658), .C1(new_n934), .C2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n733), .A2(G317), .B1(G311), .B2(new_n739), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT52), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n801), .A2(new_n514), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n393), .B1(new_n214), .B2(new_n744), .C1(new_n945), .C2(new_n754), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n741), .A2(new_n992), .B1(new_n736), .B2(new_n209), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n753), .B2(new_n724), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n733), .A2(G150), .B1(G159), .B2(new_n739), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT51), .Z(new_n1018));
  OAI22_X1  g0818(.A1(new_n801), .A2(new_n261), .B1(new_n203), .B2(new_n741), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n731), .B2(G50), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n421), .C2(new_n744), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G143), .B2(new_n759), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n297), .A3(new_n791), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n972), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n243), .A2(new_n943), .B1(new_n452), .B2(new_n224), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1025), .A2(new_n720), .A3(new_n705), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n919), .A2(new_n706), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n713), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1007), .B2(new_n939), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1008), .A2(new_n1029), .ZN(G390));
  OAI211_X1 g0830(.A(new_n891), .B(new_n611), .C1(new_n437), .C2(new_n872), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n872), .A2(new_n673), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n697), .A2(KEYINPUT88), .A3(G330), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n854), .B1(new_n1034), .B2(new_n782), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n854), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n872), .A2(new_n1036), .A3(new_n783), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n886), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n855), .B1(new_n692), .B2(new_n698), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n773), .B1(new_n668), .B2(new_n783), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n854), .B(KEYINPUT112), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n872), .B2(new_n783), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1031), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n887), .A2(new_n880), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n881), .A2(new_n1046), .A3(new_n883), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1042), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n1040), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n880), .A3(new_n850), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1039), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1037), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n782), .B1(new_n692), .B2(new_n698), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1037), .B1(new_n1055), .B2(new_n1036), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n886), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1031), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1037), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n839), .A2(new_n882), .A3(new_n849), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n882), .B1(new_n862), .B2(new_n849), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n879), .B1(new_n886), .B2(new_n854), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1050), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1060), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1054), .A2(new_n1069), .A3(new_n658), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1054), .A2(new_n1069), .A3(KEYINPUT113), .A4(new_n658), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n881), .A2(new_n703), .A3(new_n883), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n733), .A2(G128), .B1(G132), .B2(new_n739), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT114), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n745), .A2(G159), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT54), .B(G143), .Z(new_n1079));
  AOI22_X1  g0879(.A1(new_n747), .A2(new_n1079), .B1(new_n759), .B2(G125), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n297), .B1(new_n736), .B2(new_n361), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n793), .A2(G150), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT53), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G137), .C2(new_n731), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .A4(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n945), .A2(new_n209), .B1(new_n452), .B2(new_n801), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n992), .C2(new_n950), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT116), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n393), .C1(new_n203), .C2(new_n736), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G77), .A2(new_n745), .B1(new_n739), .B2(G116), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n301), .B2(new_n741), .C1(new_n514), .C2(new_n724), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1085), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n720), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1075), .A2(new_n714), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n261), .B2(new_n810), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n939), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1074), .A2(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(KEYINPUT57), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n879), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1036), .B1(new_n786), .B2(new_n773), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n863), .A2(new_n1103), .B1(new_n832), .B2(new_n639), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT117), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n407), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n387), .A2(new_n829), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1102), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1111));
  OAI21_X1  g0911(.A(G330), .B1(new_n876), .B2(new_n857), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1107), .B(new_n1108), .Z(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n884), .B2(new_n888), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1102), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n867), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1031), .B1(new_n1098), .B2(new_n1045), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1101), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1112), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1115), .A2(new_n867), .A3(new_n1116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1121), .A2(new_n1124), .A3(KEYINPUT57), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n658), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n938), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n712), .B1(new_n1114), .B2(new_n703), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n950), .A2(new_n214), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n731), .A2(G97), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n747), .A2(new_n419), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1130), .A2(new_n949), .A3(new_n998), .A4(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1129), .B(new_n1132), .C1(G283), .C2(new_n759), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G41), .B(new_n297), .C1(new_n739), .C2(G107), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n202), .C2(new_n736), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT58), .Z(new_n1136));
  OAI21_X1  g0936(.A(new_n361), .B1(new_n391), .B2(G41), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n739), .A2(G128), .ZN(new_n1138));
  INV_X1    g0938(.A(G137), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1138), .B1(new_n953), .B2(new_n744), .C1(new_n801), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n731), .A2(G132), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1079), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n741), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1140), .B(new_n1143), .C1(G125), .C2(new_n733), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT59), .ZN(new_n1145));
  AOI21_X1  g0945(.A(G33), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G41), .B1(new_n759), .B2(G124), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n268), .C2(new_n736), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n720), .B1(new_n1136), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n810), .A2(new_n361), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1128), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1127), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1126), .A2(new_n1155), .ZN(G375));
  AOI21_X1  g0956(.A(new_n713), .B1(new_n1042), .B2(new_n703), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n810), .A2(new_n203), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G128), .A2(new_n759), .B1(new_n757), .B2(G58), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n297), .C1(new_n1139), .C2(new_n740), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n733), .A2(G132), .B1(G150), .B2(new_n747), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n361), .B2(new_n744), .C1(new_n945), .C2(new_n1142), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G159), .C2(new_n793), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n733), .A2(G294), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n952), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n759), .A2(G303), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n997), .B1(G107), .B2(new_n747), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n945), .A2(new_n214), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n741), .A2(new_n452), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n393), .B1(new_n740), .B2(new_n992), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n720), .B1(new_n1163), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1157), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1058), .B2(new_n939), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1038), .A2(new_n1031), .A3(new_n1044), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1045), .A2(new_n923), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G381));
  AND2_X1   g0981(.A1(new_n1099), .A2(new_n1070), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1126), .A2(new_n1155), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1180), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n940), .A2(new_n973), .A3(new_n1029), .A4(new_n1008), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT119), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(G407));
  NAND2_X1  g0989(.A1(new_n1183), .A2(new_n640), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(G407), .A2(G213), .A3(new_n1190), .ZN(G409));
  NAND3_X1  g0991(.A1(G378), .A2(new_n1155), .A3(new_n1126), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT121), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1127), .B2(new_n1154), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n939), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT118), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1153), .B(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n923), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1121), .A2(new_n1124), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1182), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n640), .A2(G213), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT60), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1206), .A2(new_n658), .A3(new_n1060), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1176), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(G384), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n1204), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT63), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n640), .A2(G213), .A3(G2897), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1210), .B(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1192), .A2(new_n1202), .B1(G213), .B2(new_n640), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G387), .A2(G390), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(new_n1185), .ZN(new_n1222));
  XOR2_X1   g1022(.A(G393), .B(G396), .Z(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1221), .A3(new_n1185), .A4(new_n1223), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1212), .A2(KEYINPUT63), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1213), .A2(new_n1219), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  XOR2_X1   g1030(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n1217), .C2(new_n1210), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1231), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT124), .B1(new_n1211), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1203), .A2(KEYINPUT62), .A3(new_n1204), .A4(new_n1210), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1217), .A2(KEYINPUT125), .A3(KEYINPUT62), .A4(new_n1210), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1218), .B1(new_n1235), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1227), .B(KEYINPUT126), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1229), .B1(new_n1241), .B2(new_n1242), .ZN(G405));
  AOI21_X1  g1043(.A(KEYINPUT127), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1227), .B(KEYINPUT127), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G375), .A2(new_n1182), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1192), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(new_n1210), .ZN(new_n1248));
  MUX2_X1   g1048(.A(new_n1244), .B(new_n1245), .S(new_n1248), .Z(G402));
endmodule


