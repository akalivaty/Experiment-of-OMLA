//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT67), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  AND3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n209), .A2(new_n213), .B1(G1), .B2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n204), .A2(new_n205), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n214), .A2(new_n215), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n224), .B(new_n229), .C1(new_n215), .C2(new_n214), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G169), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT69), .B(G223), .Z(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n248), .A2(G1698), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G77), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n251), .A2(G222), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n264), .A3(G274), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n247), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n216), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT70), .B1(new_n275), .B2(new_n216), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n216), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n216), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G150), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n217), .A2(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n278), .B(new_n283), .C1(new_n284), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n221), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n278), .B2(new_n283), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n217), .A2(G1), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(G50), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n292), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  INV_X1    g0101(.A(new_n272), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n302), .C1(new_n262), .C2(new_n264), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n300), .B(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  OAI21_X1  g0106(.A(G200), .B1(new_n265), .B2(new_n272), .ZN(new_n307));
  OAI211_X1 g0107(.A(G190), .B(new_n302), .C1(new_n262), .C2(new_n264), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n306), .B1(new_n305), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n270), .A2(G1698), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n314), .B1(G223), .B2(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G87), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n264), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n269), .B1(new_n232), .B2(new_n271), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n318), .A3(new_n301), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(G169), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n276), .A2(new_n277), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT7), .B1(new_n255), .B2(new_n217), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n250), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G58), .A2(G68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT75), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT75), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G58), .A3(G68), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n204), .A2(new_n329), .A3(new_n331), .A4(new_n205), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n251), .B2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(KEYINPUT74), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n255), .A2(new_n340), .A3(KEYINPUT7), .A4(new_n217), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G68), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n278), .A2(new_n283), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n293), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n287), .A2(new_n297), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT76), .ZN(new_n349));
  INV_X1    g0149(.A(new_n287), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n347), .A2(new_n349), .B1(new_n293), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n321), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n336), .B2(new_n344), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT18), .B1(new_n356), .B2(new_n321), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n317), .A2(new_n318), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(G200), .B2(new_n320), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n345), .A2(new_n361), .A3(new_n352), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(KEYINPUT17), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n346), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n288), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(KEYINPUT11), .A3(new_n371), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n322), .A2(new_n294), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n297), .A2(new_n203), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT12), .B1(new_n293), .B2(G68), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(G238), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n269), .B1(new_n383), .B2(new_n271), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n232), .A2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n251), .B(new_n387), .C1(G226), .C2(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n385), .B(new_n386), .C1(new_n390), .C2(new_n264), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n264), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT13), .B1(new_n392), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n382), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n393), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n394), .A2(new_n395), .B1(new_n396), .B2(new_n301), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n394), .A2(new_n395), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n381), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(G200), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n391), .A2(G190), .A3(new_n393), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n373), .A2(new_n400), .A3(new_n380), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n251), .A2(G232), .A3(new_n258), .ZN(new_n404));
  INV_X1    g0204(.A(G107), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n251), .ZN(new_n406));
  AND2_X1   g0206(.A1(G33), .A2(G41), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n216), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n268), .A2(G274), .A3(new_n264), .ZN(new_n410));
  INV_X1    g0210(.A(new_n271), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(G244), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n247), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n350), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n288), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n322), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n375), .A2(G77), .A3(new_n298), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n294), .A2(new_n370), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n301), .A3(new_n412), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n359), .C2(new_n413), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n399), .A2(new_n402), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n313), .A2(new_n367), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G116), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n429), .A2(KEYINPUT87), .A3(G20), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT23), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n217), .B2(G107), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n405), .A2(KEYINPUT23), .A3(G20), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT87), .B1(new_n429), .B2(G20), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n251), .A2(new_n217), .A3(G87), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(KEYINPUT22), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(KEYINPUT22), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT24), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT24), .B(new_n436), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n322), .ZN(new_n444));
  INV_X1    g0244(.A(G33), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n346), .A2(G107), .A3(new_n293), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n293), .A2(G107), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT25), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n448), .A2(KEYINPUT88), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT88), .B1(new_n448), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT89), .ZN(new_n454));
  INV_X1    g0254(.A(G250), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n258), .ZN(new_n456));
  INV_X1    g0256(.A(G257), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G1698), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n458), .C1(new_n253), .C2(new_n254), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n264), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n464), .A2(G274), .A3(new_n264), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G264), .A3(new_n264), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n462), .A2(new_n463), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G169), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n471), .A2(G264), .A3(new_n264), .ZN(new_n475));
  INV_X1    g0275(.A(new_n467), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n475), .A2(new_n476), .A3(new_n461), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n474), .B1(new_n301), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT89), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n444), .B(new_n480), .C1(new_n451), .C2(new_n452), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n454), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n473), .A2(G190), .B1(G200), .B2(new_n477), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n444), .C1(new_n452), .C2(new_n451), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n293), .A2(G97), .ZN(new_n486));
  AOI211_X1 g0286(.A(new_n294), .B(new_n446), .C1(new_n278), .C2(new_n283), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(G97), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT6), .ZN(new_n489));
  AND2_X1   g0289(.A1(G97), .A2(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT6), .A2(G97), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT77), .B1(new_n493), .B2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n405), .A3(KEYINPUT6), .A4(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n324), .B2(new_n326), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n323), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT78), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI211_X1 g0302(.A(KEYINPUT78), .B(new_n323), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n488), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT81), .B(new_n488), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n471), .A2(new_n264), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n467), .B1(new_n508), .B2(new_n457), .ZN(new_n509));
  OAI211_X1 g0309(.A(G244), .B(new_n258), .C1(new_n253), .C2(new_n254), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(KEYINPUT79), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(KEYINPUT79), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n251), .A2(G244), .A3(new_n258), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n509), .B1(new_n517), .B2(new_n408), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G169), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(G179), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n506), .A2(new_n507), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n518), .A2(KEYINPUT80), .A3(G190), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT80), .B1(new_n518), .B2(G190), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G200), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n525), .A2(new_n504), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n296), .A2(G87), .A3(new_n447), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n296), .A2(KEYINPUT84), .A3(G87), .A4(new_n447), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n383), .A2(new_n258), .ZN(new_n534));
  INV_X1    g0334(.A(G244), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n536), .C1(new_n253), .C2(new_n254), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n429), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n408), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n264), .A2(G274), .A3(new_n466), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n266), .A2(G45), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(G250), .C1(new_n407), .C2(new_n216), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(new_n544), .A3(KEYINPUT82), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n264), .B1(new_n537), .B2(new_n429), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(G190), .A3(new_n548), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n251), .A2(new_n217), .A3(G68), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  INV_X1    g0353(.A(G97), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n288), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n217), .B1(new_n389), .B2(new_n553), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n491), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT83), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT83), .B1(new_n556), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n552), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n322), .B1(new_n294), .B2(new_n416), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n533), .A2(new_n550), .A3(new_n551), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n416), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n487), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n545), .A2(new_n301), .A3(new_n548), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n549), .A2(new_n247), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n522), .A2(new_n528), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n446), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n293), .B(new_n574), .C1(new_n276), .C2(new_n277), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n266), .A2(G13), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(G20), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n275), .A2(new_n216), .B1(G20), .B2(new_n573), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n515), .B(new_n217), .C1(G33), .C2(new_n554), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n575), .B1(new_n576), .B2(new_n577), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n471), .A2(G270), .A3(new_n264), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n584), .A2(new_n467), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT86), .ZN(new_n586));
  XNOR2_X1  g0386(.A(KEYINPUT85), .B(G303), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n264), .B1(new_n255), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n258), .A2(G264), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n253), .B2(new_n254), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n586), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G303), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT85), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G303), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n249), .A2(new_n594), .A3(new_n596), .A4(new_n250), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n586), .A2(new_n591), .A3(new_n597), .A4(new_n408), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n585), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n583), .A2(new_n599), .A3(new_n301), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G169), .A3(new_n582), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n599), .A2(new_n582), .A3(new_n603), .A4(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n582), .B1(new_n599), .B2(G200), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n359), .B2(new_n599), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n428), .A2(new_n485), .A3(new_n572), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n304), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT93), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT93), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n345), .A2(new_n352), .ZN(new_n614));
  INV_X1    g0414(.A(new_n321), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n354), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n399), .ZN(new_n618));
  INV_X1    g0418(.A(new_n423), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n402), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n611), .B(new_n617), .C1(new_n620), .C2(new_n366), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n305), .A2(new_n309), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n610), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n547), .A2(new_n543), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n247), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n566), .A2(new_n567), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n563), .A2(new_n569), .ZN(new_n632));
  XNOR2_X1  g0432(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n522), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(G200), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n533), .A2(new_n551), .A3(new_n562), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n520), .A2(new_n521), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n504), .A4(new_n630), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n522), .A2(new_n528), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n453), .A2(new_n479), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n605), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT91), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n484), .A2(new_n630), .A3(new_n637), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n644), .A2(new_n648), .A3(new_n605), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n643), .A2(new_n646), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n626), .B1(new_n428), .B2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(new_n605), .ZN(new_n653));
  OR3_X1    g0453(.A1(new_n576), .A2(KEYINPUT27), .A3(G20), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT27), .B1(new_n576), .B2(G20), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g0456(.A(KEYINPUT94), .B(G343), .Z(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n583), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT95), .B1(new_n653), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n608), .B2(new_n660), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n653), .A2(KEYINPUT95), .A3(new_n660), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n482), .A2(new_n659), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n482), .A2(new_n484), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n454), .A2(new_n481), .A3(new_n658), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n653), .A2(new_n659), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n485), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n453), .A2(new_n479), .A3(new_n659), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n226), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n558), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n223), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n498), .A2(new_n499), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n322), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT78), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n500), .A2(new_n501), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT81), .B1(new_n690), .B2(new_n488), .ZN(new_n691));
  INV_X1    g0491(.A(new_n507), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n638), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n633), .B1(new_n693), .B2(new_n570), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n637), .A2(new_n630), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n638), .A2(new_n504), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(KEYINPUT26), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n631), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT96), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n522), .B2(new_n528), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n523), .A2(new_n524), .ZN(new_n701));
  INV_X1    g0501(.A(new_n527), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n690), .A3(new_n488), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n693), .A2(KEYINPUT96), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n482), .A2(new_n605), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n700), .A2(new_n704), .A3(new_n647), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n658), .B1(new_n698), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n658), .B1(new_n642), .B2(new_n650), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n584), .A2(new_n467), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n591), .A2(new_n597), .A3(new_n408), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT86), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n588), .A2(new_n586), .A3(new_n591), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n475), .A2(new_n461), .A3(new_n301), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n548), .A3(new_n545), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n712), .B1(new_n719), .B2(new_n519), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT82), .B1(new_n539), .B2(new_n544), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n547), .A2(new_n543), .A3(new_n546), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G250), .A2(G1698), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n457), .B2(G1698), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n724), .A2(new_n251), .B1(G33), .B2(G294), .ZN(new_n725));
  OAI211_X1 g0525(.A(G179), .B(new_n472), .C1(new_n725), .C2(new_n264), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n721), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .A3(new_n518), .A4(new_n717), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n477), .A2(G179), .A3(new_n627), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n519), .A3(new_n599), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n720), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n658), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n602), .A2(new_n604), .ZN(new_n736));
  INV_X1    g0536(.A(new_n600), .ZN(new_n737));
  AND4_X1   g0537(.A1(new_n736), .A2(new_n737), .A3(new_n607), .A4(new_n659), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n693), .A2(new_n738), .A3(new_n703), .A4(new_n632), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n734), .B(new_n735), .C1(new_n739), .C2(new_n485), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n709), .A2(new_n711), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n685), .B1(new_n743), .B2(G1), .ZN(G364));
  NAND2_X1  g0544(.A1(new_n217), .A2(G13), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT98), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n266), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n665), .B1(new_n680), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n664), .A2(G330), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n664), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n216), .B1(G20), .B2(new_n247), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n679), .A2(new_n251), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n242), .A2(new_n465), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT99), .Z(new_n761));
  AOI211_X1 g0561(.A(new_n759), .B(new_n761), .C1(new_n465), .C2(new_n222), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n251), .A2(new_n226), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n226), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n757), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n217), .A2(G179), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT32), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(new_n359), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n217), .A2(new_n301), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n773), .B1(new_n405), .B2(new_n774), .C1(new_n203), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(new_n768), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n775), .A2(G190), .A3(new_n526), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n251), .B1(new_n780), .B2(new_n370), .C1(new_n202), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(new_n359), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n359), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n217), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n221), .B1(new_n554), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n772), .A2(KEYINPUT32), .B1(new_n557), .B2(new_n788), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n779), .A2(new_n782), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G317), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT33), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(KEYINPUT33), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n777), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n795), .B2(new_n786), .C1(new_n593), .C2(new_n788), .ZN(new_n796));
  INV_X1    g0596(.A(new_n781), .ZN(new_n797));
  INV_X1    g0597(.A(new_n769), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G322), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n255), .C1(new_n800), .C2(new_n780), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(G326), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n774), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n796), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n790), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT100), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT100), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n807), .A2(new_n808), .A3(new_n756), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n748), .A2(new_n680), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n766), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n749), .A2(new_n750), .B1(new_n755), .B2(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n421), .A2(new_n658), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n426), .A2(new_n423), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT102), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT102), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n426), .A2(new_n816), .A3(new_n423), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n658), .B(new_n819), .C1(new_n642), .C2(new_n650), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n619), .A2(new_n658), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n815), .A2(new_n822), .A3(new_n817), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT103), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n710), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n810), .B1(new_n825), .B2(new_n741), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n741), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n756), .A2(new_n751), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n810), .B1(G77), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n784), .A2(new_n593), .B1(new_n788), .B2(new_n405), .ZN(new_n831));
  INV_X1    g0631(.A(new_n774), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(G87), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n251), .B1(new_n797), .B2(G294), .ZN(new_n834));
  INV_X1    g0634(.A(new_n780), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G116), .A2(new_n835), .B1(new_n798), .B2(G311), .ZN(new_n836));
  INV_X1    g0636(.A(new_n786), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G97), .A2(new_n837), .B1(new_n777), .B2(G283), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n833), .A2(new_n834), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n797), .A2(G143), .B1(new_n835), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n778), .B2(new_n841), .C1(new_n842), .C2(new_n784), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n251), .B1(new_n769), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G68), .B2(new_n832), .ZN(new_n848));
  INV_X1    g0648(.A(new_n788), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n837), .A2(G58), .B1(new_n849), .B2(G50), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n843), .A2(new_n844), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n839), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n830), .B1(new_n853), .B2(new_n756), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n823), .B2(new_n752), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n827), .A2(new_n855), .ZN(G384));
  AND2_X1   g0656(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(new_n573), .A4(new_n219), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n222), .A2(G77), .A3(new_n331), .A4(new_n329), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n221), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n266), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n709), .A2(new_n711), .ZN(new_n865));
  INV_X1    g0665(.A(new_n428), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n626), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(new_n366), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n617), .A2(new_n870), .A3(new_n611), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n656), .B1(new_n345), .B2(new_n352), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n345), .A2(new_n361), .A3(new_n352), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(new_n353), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n362), .B(KEYINPUT93), .C1(new_n356), .C2(new_n656), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(KEYINPUT37), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n362), .B1(new_n356), .B2(new_n656), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NOR4_X1   g0680(.A1(new_n879), .A2(KEYINPUT93), .A3(new_n880), .A4(new_n353), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n332), .A2(G20), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n285), .A2(G159), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(G68), .B2(new_n342), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n346), .B1(new_n887), .B2(KEYINPUT16), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n343), .A2(new_n333), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n335), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n351), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n362), .B1(new_n891), .B2(new_n321), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n656), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n875), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n893), .B1(new_n358), .B2(new_n366), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n869), .B1(new_n883), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n618), .A2(new_n659), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n381), .A2(new_n658), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n399), .A2(new_n402), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n381), .B(new_n658), .C1(new_n397), .C2(new_n398), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n423), .A2(new_n658), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n908), .B(new_n912), .C1(new_n820), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n617), .A2(new_n611), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n656), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n907), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n868), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(G330), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(new_n823), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT31), .B1(new_n731), .B2(new_n658), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(KEYINPUT104), .B2(new_n735), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n733), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n667), .A2(new_n571), .A3(new_n738), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(KEYINPUT40), .C1(new_n883), .C2(new_n899), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n734), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n923), .C1(new_n485), .C2(new_n739), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n912), .A2(new_n823), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n899), .C2(new_n904), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n931), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n428), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n919), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n918), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n266), .B2(new_n746), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n918), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n864), .B1(new_n943), .B2(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n533), .A2(new_n562), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n658), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n695), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT105), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT105), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(new_n630), .C2(new_n947), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(new_n754), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n757), .B1(new_n226), .B2(new_n416), .C1(new_n238), .C2(new_n759), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n810), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n781), .A2(new_n841), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n786), .A2(new_n203), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(G143), .C2(new_n783), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(KEYINPUT109), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(KEYINPUT109), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n251), .B1(new_n769), .B2(new_n842), .C1(new_n221), .C2(new_n780), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n832), .A2(G77), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n202), .B2(new_n788), .C1(new_n778), .C2(new_n770), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n587), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n797), .A2(new_n964), .B1(new_n798), .B2(G317), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n849), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n251), .B1(new_n835), .B2(G283), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n778), .A2(new_n795), .B1(new_n774), .B2(new_n554), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n784), .A2(new_n800), .B1(new_n405), .B2(new_n786), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n849), .B2(G116), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  AOI21_X1  g0774(.A(new_n954), .B1(new_n974), .B2(new_n756), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n952), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n504), .A2(new_n658), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n700), .A2(new_n704), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n696), .A2(new_n658), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n671), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n693), .B1(new_n984), .B2(new_n482), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n659), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n984), .B2(new_n674), .ZN(new_n989));
  OAI211_X1 g0789(.A(KEYINPUT42), .B(new_n673), .C1(new_n982), .C2(new_n983), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n987), .A2(new_n991), .A3(KEYINPUT107), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n987), .A2(new_n991), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n951), .B(KEYINPUT43), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n985), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n985), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n978), .A2(new_n980), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT106), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n676), .A3(new_n981), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n984), .B2(new_n676), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n677), .B(KEYINPUT45), .C1(new_n982), .C2(new_n983), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n670), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n669), .A2(new_n672), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n674), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n665), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1009), .A2(new_n1013), .A3(new_n671), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1015), .A2(new_n743), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n743), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n680), .B(KEYINPUT41), .Z(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n748), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1004), .A2(new_n1025), .A3(KEYINPUT108), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT108), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n747), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n997), .A2(new_n985), .A3(new_n1000), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n1001), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n976), .B1(new_n1026), .B2(new_n1032), .ZN(G387));
  AND2_X1   g0833(.A1(new_n743), .A2(new_n1019), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n681), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n743), .B2(new_n1019), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n669), .A2(new_n753), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n763), .A2(new_n682), .B1(G107), .B2(new_n226), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n235), .A2(new_n465), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n682), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G45), .B(new_n1040), .C1(G68), .C2(G77), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n287), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n759), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1038), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n757), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n810), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT110), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n780), .A2(new_n203), .B1(new_n769), .B2(new_n841), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n255), .B(new_n1049), .C1(G50), .C2(new_n797), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n849), .A2(G77), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n564), .A2(new_n837), .B1(new_n777), .B2(new_n350), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n783), .A2(G159), .B1(new_n832), .B2(G97), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n797), .A2(G317), .B1(new_n835), .B2(new_n964), .ZN(new_n1055));
  INV_X1    g0855(.A(G322), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n784), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G311), .B2(new_n777), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n786), .A2(new_n803), .B1(new_n788), .B2(new_n795), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT111), .Z(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n251), .B1(new_n798), .B2(G326), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n573), .C2(new_n774), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1054), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1048), .B1(new_n1070), .B2(new_n756), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1019), .A2(new_n748), .B1(new_n1037), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1036), .A2(new_n1072), .ZN(G393));
  AND2_X1   g0873(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n748), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n982), .A2(new_n754), .A3(new_n983), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n245), .A2(new_n758), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n757), .C1(new_n554), .C2(new_n226), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n784), .A2(new_n841), .B1(new_n770), .B2(new_n781), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n778), .A2(new_n221), .B1(new_n774), .B2(new_n557), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n255), .B1(new_n798), .B2(G143), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n287), .B2(new_n780), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n786), .A2(new_n370), .B1(new_n788), .B2(new_n203), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n784), .A2(new_n791), .B1(new_n800), .B2(new_n781), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n778), .A2(new_n587), .B1(new_n573), .B2(new_n786), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n255), .B1(new_n769), .B2(new_n1056), .C1(new_n795), .C2(new_n780), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n405), .A2(new_n774), .B1(new_n788), .B2(new_n803), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1080), .A2(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n756), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n810), .B(new_n1078), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT114), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1075), .B1(new_n1076), .B2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1074), .A2(new_n1034), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1021), .A2(new_n680), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  INV_X1    g0901(.A(KEYINPUT115), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n937), .A2(new_n919), .A3(new_n920), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n912), .B1(new_n820), .B2(new_n913), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1104), .A2(new_n901), .B1(new_n900), .B2(new_n906), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n901), .B1(new_n883), .B2(new_n899), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n707), .A2(new_n818), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n913), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1109), .B2(new_n912), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1102), .B(new_n1103), .C1(new_n1105), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n913), .B1(new_n710), .B2(new_n818), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n912), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n901), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n900), .A2(new_n906), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n883), .A2(new_n899), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n913), .B1(new_n707), .B2(new_n818), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n901), .B(new_n1117), .C1(new_n1118), .C2(new_n1113), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n740), .A2(G330), .A3(new_n823), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1116), .B(new_n1119), .C1(new_n1113), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1102), .B1(new_n1123), .B2(new_n1103), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n824), .A2(G330), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n912), .B1(new_n1126), .B2(new_n931), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1120), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n912), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n927), .A2(G330), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1128), .B2(new_n912), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1112), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1129), .A2(new_n1118), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n938), .A2(G330), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT116), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n626), .A3(new_n867), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n680), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n781), .A2(new_n846), .B1(new_n780), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n255), .B(new_n1143), .C1(G125), .C2(new_n798), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n788), .A2(new_n841), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n777), .A2(G137), .B1(new_n832), .B2(G50), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n786), .A2(new_n770), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G128), .B2(new_n783), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n786), .A2(new_n370), .B1(new_n781), .B2(new_n573), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n255), .B1(new_n780), .B2(new_n554), .C1(new_n557), .C2(new_n788), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n405), .A2(new_n778), .B1(new_n784), .B2(new_n803), .ZN(new_n1154));
  OR3_X1    g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n774), .A2(new_n203), .B1(new_n769), .B2(new_n795), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT117), .Z(new_n1157));
  OAI21_X1  g0957(.A(new_n1150), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n756), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n810), .C1(new_n350), .C2(new_n829), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1115), .B2(new_n751), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1125), .B2(new_n748), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1141), .A2(new_n1162), .ZN(G378));
  NAND3_X1  g0963(.A1(new_n928), .A2(new_n935), .A3(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n656), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n300), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT119), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n625), .B2(new_n304), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n304), .B(new_n1171), .C1(new_n310), .C2(new_n311), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1168), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1171), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n312), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1167), .A3(new_n1173), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n928), .A2(new_n935), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1166), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AND4_X1   g0982(.A1(G330), .A2(new_n928), .A3(new_n935), .A4(new_n1179), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n917), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n917), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1182), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1186), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT122), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1186), .B(KEYINPUT122), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1137), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1140), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1186), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1137), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n680), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1180), .A2(new_n751), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n810), .B1(G50), .B2(new_n829), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n784), .A2(new_n573), .B1(new_n774), .B2(new_n202), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G97), .B2(new_n777), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n251), .A2(G41), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G283), .B2(new_n798), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n797), .A2(G107), .B1(new_n835), .B2(new_n564), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n956), .B1(G77), .B2(new_n849), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1209), .B(new_n221), .C1(G33), .C2(G41), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n783), .A2(G125), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n778), .B2(new_n846), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n797), .A2(G128), .B1(new_n835), .B2(G137), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n788), .B2(new_n1142), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G150), .C2(new_n837), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n832), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1217), .B1(new_n1214), .B2(new_n1213), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1206), .B1(new_n1229), .B2(new_n756), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1205), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1195), .B2(new_n748), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1204), .A2(new_n1233), .ZN(G375));
  INV_X1    g1034(.A(new_n1138), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1024), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n810), .B1(G68), .B2(new_n829), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n573), .A2(new_n778), .B1(new_n784), .B2(new_n795), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G97), .B2(new_n849), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n837), .A2(new_n564), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n781), .A2(new_n803), .B1(new_n780), .B2(new_n405), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n251), .B(new_n1242), .C1(G303), .C2(new_n798), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n961), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n255), .B1(new_n798), .B2(G128), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n842), .B2(new_n781), .C1(new_n841), .C2(new_n780), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n778), .A2(new_n1142), .B1(new_n774), .B2(new_n202), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G50), .A2(new_n837), .B1(new_n783), .B2(G132), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n770), .C2(new_n788), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1093), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(new_n1250), .A3(KEYINPUT123), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1238), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n912), .B2(new_n752), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1133), .B2(new_n747), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(new_n1258), .ZN(G381));
  NOR2_X1   g1059(.A1(G393), .A2(G396), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G381), .A2(G384), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1100), .A3(new_n1261), .ZN(new_n1262));
  OR4_X1    g1062(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1262), .ZN(G407));
  AND2_X1   g1063(.A1(new_n1141), .A2(new_n1162), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n657), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G375), .C2(new_n1267), .ZN(G409));
  XOR2_X1   g1068(.A(G393), .B(G396), .Z(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n976), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT108), .B1(new_n1004), .B2(new_n1025), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1029), .A2(new_n1031), .A3(new_n1027), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1271), .B(new_n1100), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n1275), .B2(new_n976), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(new_n1100), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n976), .A3(G390), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1269), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1233), .C1(new_n1198), .C2(new_n1203), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1023), .B(new_n1202), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1200), .A2(new_n748), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1231), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1264), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1266), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n681), .B(new_n1138), .C1(new_n1289), .C2(new_n1236), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1133), .A2(new_n1137), .A3(KEYINPUT60), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT125), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1257), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  XOR2_X1   g1096(.A(G384), .B(KEYINPUT126), .Z(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1282), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1283), .A2(new_n1287), .A3(KEYINPUT124), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1265), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1266), .A2(G2897), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1296), .B(new_n1307), .C1(new_n1293), .C2(new_n1297), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(G2897), .A3(new_n1266), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1304), .A2(new_n1265), .A3(new_n1299), .A4(new_n1305), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1301), .A2(new_n1310), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1308), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1281), .B1(new_n1315), .B2(new_n1288), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1311), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1288), .A2(KEYINPUT62), .A3(new_n1299), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1316), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1314), .B1(new_n1320), .B2(new_n1321), .ZN(G405));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G378), .B1(new_n1204), .B2(new_n1233), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1283), .ZN(new_n1326));
  OR3_X1    g1126(.A1(new_n1325), .A2(new_n1299), .A3(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1299), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT127), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1324), .A2(new_n1327), .A3(new_n1328), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(KEYINPUT127), .A3(new_n1329), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(G402));
endmodule


