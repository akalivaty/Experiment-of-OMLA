//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n538, new_n539, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT68), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT68), .B1(new_n466), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n473), .B2(G2105), .ZN(G160));
  NAND2_X1  g049(.A1(new_n461), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n461), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n489), .B2(new_n478), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n478), .C1(new_n469), .C2(new_n470), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n501), .A2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  AOI22_X1  g086(.A1(new_n504), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(new_n497), .ZN(new_n513));
  INV_X1    g088(.A(new_n507), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(G51), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XOR2_X1   g091(.A(new_n516), .B(KEYINPUT7), .Z(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(G286));
  INV_X1    g094(.A(G286), .ZN(G168));
  AOI22_X1  g095(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n500), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G90), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n505), .A2(new_n523), .B1(new_n507), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G171));
  NAND2_X1  g101(.A1(G68), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G56), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n497), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT70), .ZN(new_n531));
  INV_X1    g106(.A(new_n505), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G81), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n514), .A2(G43), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n538), .A2(new_n542), .ZN(G188));
  XNOR2_X1  g118(.A(new_n497), .B(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G65), .ZN(new_n545));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n500), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n548));
  NAND3_X1  g123(.A1(new_n514), .A2(G53), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n532), .A2(G91), .ZN(new_n550));
  NOR2_X1   g125(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n507), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  NAND2_X1  g132(.A1(new_n532), .A2(G87), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n514), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  OAI211_X1 g136(.A(G48), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  AOI22_X1  g140(.A1(G86), .A2(new_n532), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n497), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT75), .ZN(G305));
  AOI22_X1  g147(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n500), .ZN(new_n574));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n505), .A2(new_n575), .B1(new_n507), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G290));
  INV_X1    g154(.A(G868), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(G171), .B2(new_n580), .ZN(new_n581));
  OR3_X1    g156(.A1(G171), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n532), .A2(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  NAND2_X1  g159(.A1(new_n514), .A2(G54), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n544), .A2(G66), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT77), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n581), .B(new_n582), .C1(new_n590), .C2(G868), .ZN(G284));
  OAI211_X1 g166(.A(new_n581), .B(new_n582), .C1(new_n590), .C2(G868), .ZN(G321));
  NAND2_X1  g167(.A1(G286), .A2(G868), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n555), .B(KEYINPUT78), .Z(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(G868), .ZN(G297));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(G868), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n536), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g177(.A(KEYINPUT68), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n467), .A2(G2104), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT68), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n465), .A2(G2105), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n476), .A2(G123), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT79), .ZN(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n480), .A2(G135), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XOR2_X1   g199(.A(G2443), .B(G2446), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n628), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  OAI21_X1  g215(.A(KEYINPUT17), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n640), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n642), .A2(new_n638), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n637), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n644), .B(new_n645), .C1(new_n643), .C2(new_n637), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(new_n613), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT81), .B(G2096), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT82), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n652), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(G1981), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1991), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n667), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n678), .A3(new_n676), .ZN(new_n681));
  AND2_X1   g256(.A1(KEYINPUT87), .A2(G16), .ZN(new_n682));
  NOR2_X1   g257(.A1(KEYINPUT87), .A2(G16), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G166), .B2(new_n685), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT33), .Z(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G1976), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(G1976), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n687), .A2(G1971), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n680), .A2(new_n681), .A3(new_n688), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G119), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n480), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(new_n478), .B2(G107), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT85), .B(G29), .ZN(new_n706));
  MUX2_X1   g281(.A(G25), .B(new_n705), .S(new_n706), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n685), .A2(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n578), .B2(new_n685), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n710), .B1(new_n712), .B2(G1986), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G1986), .B2(new_n712), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n698), .B2(KEYINPUT34), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n699), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n536), .A2(new_n685), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G19), .B2(new_n685), .ZN(new_n720));
  INV_X1    g295(.A(G1341), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n699), .A2(new_n715), .A3(KEYINPUT36), .A4(new_n709), .ZN(new_n723));
  NOR3_X1   g298(.A1(KEYINPUT90), .A2(G29), .A3(G33), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n608), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT92), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT92), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(G2105), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n609), .A2(G103), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  INV_X1    g307(.A(G139), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n479), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n724), .B1(new_n737), .B2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(KEYINPUT90), .B1(G29), .B2(G33), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(G2072), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT95), .Z(new_n741));
  AOI21_X1  g316(.A(G2072), .B1(new_n738), .B2(new_n739), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G168), .B2(G16), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G1966), .ZN(new_n746));
  NOR2_X1   g321(.A1(G5), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G171), .B2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(G1961), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n620), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT30), .B(G28), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n706), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(G129), .A2(new_n476), .B1(new_n480), .B2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n609), .A2(G105), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G32), .B(new_n758), .S(G29), .Z(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  OAI211_X1 g335(.A(new_n749), .B(new_n753), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n476), .A2(G128), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n480), .A2(G140), .ZN(new_n763));
  NOR2_X1   g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G26), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n706), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(G29), .B1(KEYINPUT28), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT28), .B2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n761), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  MUX2_X1   g348(.A(G35), .B(new_n484), .S(new_n706), .Z(new_n774));
  XOR2_X1   g349(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n745), .A2(G1966), .B1(new_n759), .B2(new_n760), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G1961), .ZN(new_n781));
  INV_X1    g356(.A(new_n748), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n685), .A2(KEYINPUT23), .A3(G20), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G20), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n684), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n555), .C2(new_n689), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT98), .B(G1956), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT99), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n772), .A2(new_n773), .A3(new_n783), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(G160), .A2(G29), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT24), .B(G34), .Z(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n706), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n590), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G1348), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n721), .B2(new_n720), .ZN(new_n803));
  INV_X1    g378(.A(G27), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n706), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n486), .A2(new_n487), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n478), .ZN(new_n807));
  INV_X1    g382(.A(G138), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n808), .B(G2105), .C1(new_n606), .C2(new_n607), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT4), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n811));
  NAND2_X1  g386(.A1(G114), .A2(G2104), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n807), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n805), .B1(new_n815), .B2(new_n706), .ZN(new_n816));
  MUX2_X1   g391(.A(new_n805), .B(new_n816), .S(KEYINPUT96), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G2078), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n776), .A2(new_n777), .B1(new_n796), .B2(new_n795), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n801), .B2(new_n800), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n803), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n741), .A2(new_n743), .A3(new_n792), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n718), .A2(new_n722), .A3(new_n723), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  AOI22_X1  g399(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n500), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n505), .A2(new_n827), .B1(new_n507), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n590), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n536), .A2(new_n831), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n535), .A2(new_n830), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT39), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n835), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(G860), .ZN(G145));
  XNOR2_X1  g416(.A(G162), .B(G160), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n736), .B(new_n705), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n611), .B(KEYINPUT100), .ZN(new_n844));
  XNOR2_X1  g419(.A(G164), .B(new_n766), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n844), .B(new_n845), .Z(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n737), .A2(new_n705), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n730), .A2(new_n705), .A3(new_n735), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n476), .A2(G130), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n480), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n758), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n848), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n848), .B2(new_n851), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n859), .A2(new_n860), .A3(new_n620), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n843), .A2(new_n847), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n849), .A2(new_n846), .A3(new_n850), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n848), .A2(new_n851), .A3(new_n858), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n750), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n842), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n620), .B1(new_n859), .B2(new_n860), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n750), .A3(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(new_n842), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT40), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n867), .A2(new_n875), .A3(new_n868), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G395));
  NAND2_X1  g452(.A1(new_n590), .A2(new_n555), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT41), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n599), .B(new_n838), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n883), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n885), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n691), .B(G303), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G305), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(new_n578), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n578), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT42), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n888), .A3(new_n887), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n580), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n830), .A2(G868), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n901), .A2(KEYINPUT102), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT102), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  OR2_X1    g480(.A1(new_n901), .A2(new_n902), .ZN(G331));
  NAND3_X1  g481(.A1(new_n836), .A2(G301), .A3(new_n837), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G301), .B1(new_n836), .B2(new_n837), .ZN(new_n909));
  OAI21_X1  g484(.A(G286), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(G168), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n882), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n910), .A2(new_n912), .A3(new_n880), .A4(new_n878), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n893), .A3(new_n892), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n894), .A3(new_n915), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n868), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  XOR2_X1   g495(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n917), .A2(new_n868), .A3(new_n922), .A4(new_n918), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(KEYINPUT44), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n921), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n923), .ZN(new_n926));
  XOR2_X1   g501(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G397));
  XOR2_X1   g503(.A(KEYINPUT105), .B(G1384), .Z(new_n929));
  AOI21_X1  g504(.A(new_n478), .B1(new_n811), .B2(new_n812), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n491), .B1(new_n810), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n931), .B2(new_n807), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n478), .B1(new_n471), .B2(new_n472), .ZN(new_n938));
  INV_X1    g513(.A(G40), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(new_n464), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(G1996), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT127), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n942), .B(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n941), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n766), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n758), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n945), .B(new_n950), .C1(new_n943), .C2(KEYINPUT46), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  NOR2_X1   g527(.A1(new_n766), .A2(G2067), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n949), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n758), .B(G1996), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n955), .A2(new_n956), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n705), .A2(new_n708), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n705), .A2(new_n708), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n946), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1986), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n578), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT107), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n941), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT48), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n960), .A2(new_n941), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n952), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n691), .A2(G1976), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND4_X1  g548(.A1(G160), .A2(new_n815), .A3(G40), .A4(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(KEYINPUT112), .A3(G8), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT112), .B1(new_n974), .B2(G8), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT113), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n972), .B(new_n979), .C1(new_n975), .C2(new_n976), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  NAND3_X1  g558(.A1(G288), .A2(new_n978), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n532), .A2(G86), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n564), .A2(new_n565), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n664), .A4(new_n570), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n566), .A2(KEYINPUT114), .A3(new_n664), .A4(new_n570), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n571), .A2(G1981), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n995), .A2(new_n996), .B1(new_n975), .B2(new_n976), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n929), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n815), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n932), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n464), .ZN(new_n1005));
  INV_X1    g580(.A(new_n472), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n608), .B2(G125), .ZN(new_n1007));
  OAI211_X1 g582(.A(G40), .B(new_n1005), .C1(new_n1007), .C2(new_n478), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n815), .A2(new_n973), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n934), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1971), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n931), .B2(new_n807), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n777), .A3(new_n1015), .A4(new_n940), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT55), .Z(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n934), .B1(G164), .B2(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n940), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1021), .B(new_n1016), .C1(new_n1024), .C2(G1971), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1018), .A2(G8), .A3(new_n1020), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1020), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1030));
  INV_X1    g605(.A(G2078), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1022), .A4(new_n940), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT123), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1010), .A2(new_n1034), .A3(new_n1031), .A4(new_n1030), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1035), .A3(KEYINPUT53), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1014), .A2(new_n940), .A3(new_n1015), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n781), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT110), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n1039));
  NOR4_X1   g614(.A1(G164), .A2(new_n1001), .A3(new_n934), .A4(new_n929), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1010), .B(new_n1031), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G171), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n998), .A2(new_n1026), .A3(new_n1029), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1010), .A2(new_n1030), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n796), .A2(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n1051), .B2(G168), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1051), .B2(G168), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1048), .A2(new_n796), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(G168), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1055), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n971), .B1(new_n1047), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1026), .A2(new_n997), .A3(new_n1029), .A4(new_n985), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1055), .A2(new_n1061), .A3(new_n1056), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(KEYINPUT126), .A3(new_n1068), .A4(new_n1046), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1010), .B(new_n1071), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1037), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  INV_X1    g650(.A(new_n547), .ZN(new_n1076));
  INV_X1    g651(.A(new_n554), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n547), .A2(new_n554), .A3(KEYINPUT57), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1072), .A2(new_n1074), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(KEYINPUT119), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(KEYINPUT119), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1037), .A2(new_n801), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n974), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n940), .A2(new_n1012), .A3(KEYINPUT118), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n947), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n879), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1081), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1010), .B(new_n666), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NOR4_X1   g669(.A1(new_n1008), .A2(G164), .A3(new_n1087), .A4(G1384), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT118), .B1(new_n940), .B2(new_n1012), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT59), .B1(new_n1098), .B2(new_n536), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1100), .B(new_n535), .C1(new_n1093), .C2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  AND4_X1   g677(.A1(new_n1102), .A2(new_n1086), .A3(new_n1090), .A4(new_n590), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1072), .A2(new_n1080), .A3(new_n1074), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1080), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1086), .A2(new_n1090), .A3(new_n879), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT60), .B1(new_n1111), .B2(new_n1091), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT120), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1104), .A2(new_n1110), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1081), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1072), .A2(new_n1074), .A3(new_n1080), .A4(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT122), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n1120), .A3(KEYINPUT61), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1092), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1066), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1124));
  AOI21_X1  g699(.A(G2078), .B1(new_n940), .B2(KEYINPUT124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1042), .B1(new_n1008), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n936), .A2(new_n1004), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(new_n1043), .A3(G301), .A4(new_n1038), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n1045), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1043), .A3(new_n1038), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1036), .A2(new_n1043), .A3(G301), .A4(new_n1038), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT54), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT125), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1136), .A3(KEYINPUT54), .A4(new_n1133), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1130), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1123), .A2(new_n1124), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1070), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1018), .A2(G8), .A3(new_n1025), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1028), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1059), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1026), .A2(new_n997), .A3(new_n985), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT116), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1054), .A2(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1066), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1143), .B1(new_n1141), .B2(new_n1028), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n998), .A4(new_n1026), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n997), .A2(new_n983), .A3(new_n691), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n992), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT115), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n975), .A2(new_n976), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1026), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1158), .A2(new_n1159), .B1(new_n1160), .B2(new_n998), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT117), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1154), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1140), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n966), .B1(new_n964), .B2(new_n578), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n946), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n958), .A2(new_n962), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT109), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n970), .B1(new_n1166), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g746(.A(G401), .B1(new_n925), .B2(new_n923), .ZN(new_n1173));
  NOR3_X1   g747(.A1(G229), .A2(new_n459), .A3(G227), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n1173), .A2(new_n873), .A3(new_n1174), .ZN(G308));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n873), .A3(new_n1174), .ZN(G225));
endmodule


