//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT74), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT70), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(new_n207), .B2(G120gat), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT71), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G127gat), .ZN(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G134gat), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n221), .B(new_n208), .C1(new_n210), .C2(new_n212), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n214), .A2(new_n220), .A3(KEYINPUT73), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n214), .A2(new_n222), .A3(new_n220), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G127gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G127gat), .B2(new_n216), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n212), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n211), .A2(G113gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT1), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(new_n229), .B2(new_n230), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n223), .A2(new_n226), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n245));
  NOR2_X1   g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT23), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(KEYINPUT23), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n243), .A2(new_n249), .A3(KEYINPUT25), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(new_n244), .ZN(new_n253));
  INV_X1    g052(.A(G169gat), .ZN(new_n254));
  INV_X1    g053(.A(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n246), .A2(new_n259), .A3(KEYINPUT23), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n250), .A2(KEYINPUT64), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n252), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT27), .B(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n268), .B2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n270), .C1(KEYINPUT67), .C2(KEYINPUT28), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n256), .A2(KEYINPUT26), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n244), .B1(new_n246), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n241), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n265), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n236), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n226), .A2(new_n223), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n231), .A2(new_n235), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n276), .B1(new_n269), .B2(new_n271), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n251), .B2(new_n264), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G227gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n206), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n278), .A2(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(new_n287), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT34), .B(new_n287), .C1(new_n278), .C2(new_n284), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n288), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n300));
  INV_X1    g099(.A(new_n298), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n299), .A2(KEYINPUT36), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT36), .B1(new_n299), .B2(new_n302), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT0), .ZN(new_n307));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n313));
  XNOR2_X1  g112(.A(G155gat), .B(G162gat), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  OR3_X1    g114(.A1(new_n315), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT80), .B(G162gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(G155gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n314), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(KEYINPUT2), .B2(new_n312), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n281), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n321), .A2(new_n323), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n279), .A3(new_n280), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n329), .B(KEYINPUT82), .Z(new_n330));
  AOI21_X1  g129(.A(new_n311), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n323), .C1(new_n317), .C2(new_n320), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT81), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n281), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n326), .ZN(new_n339));
  INV_X1    g138(.A(new_n330), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n336), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n331), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n311), .A3(new_n340), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n337), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT4), .B1(new_n236), .B2(new_n326), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT83), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(new_n347), .A3(new_n339), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n343), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n310), .B1(new_n342), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(new_n348), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n338), .B2(new_n339), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n341), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n309), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(KEYINPUT6), .B(new_n310), .C1(new_n342), .C2(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n360), .B(KEYINPUT76), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n283), .B2(KEYINPUT29), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n283), .B2(new_n360), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G197gat), .B(G204gat), .Z(new_n369));
  AOI21_X1  g168(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n373), .B(KEYINPUT75), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n360), .B1(new_n283), .B2(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n277), .A2(new_n363), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  AND3_X1   g181(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n382), .A2(KEYINPUT38), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n378), .A2(new_n377), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n375), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n374), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n385), .A3(new_n379), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n359), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT88), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n379), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT37), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396));
  INV_X1    g195(.A(new_n382), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n385), .B1(new_n376), .B2(new_n379), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT89), .B1(new_n399), .B2(new_n382), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n390), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n358), .A2(new_n405), .A3(new_n359), .A4(new_n391), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(KEYINPUT90), .A3(KEYINPUT38), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n393), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT85), .B1(G228gat), .B2(G233gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n332), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n324), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n334), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n413), .B2(new_n374), .ZN(new_n414));
  NAND3_X1  g213(.A1(KEYINPUT85), .A2(G228gat), .A3(G233gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G22gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n414), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n417), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n417), .A2(new_n422), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT39), .B1(new_n328), .B2(new_n330), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT87), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(KEYINPUT39), .C1(new_n328), .C2(new_n330), .ZN(new_n430));
  INV_X1    g229(.A(new_n336), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n346), .B2(new_n348), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n428), .B(new_n430), .C1(new_n432), .C2(new_n340), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n336), .B1(new_n352), .B2(new_n353), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n330), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT40), .A4(new_n309), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n382), .B1(new_n376), .B2(new_n379), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n383), .B2(KEYINPUT30), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT78), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n437), .A2(new_n445), .A3(new_n350), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n433), .A2(new_n436), .A3(new_n309), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n426), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n305), .B1(new_n408), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n358), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT84), .B1(new_n358), .B2(new_n359), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n426), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n299), .A2(new_n302), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n426), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n358), .A2(new_n359), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n452), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n445), .B1(new_n465), .B2(new_n453), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n426), .A2(new_n459), .A3(new_n463), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n462), .A2(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(KEYINPUT91), .A3(new_n468), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G113gat), .B(G141gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(G197gat), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT11), .B(G169gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n477), .B(KEYINPUT12), .Z(new_n478));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n480));
  INV_X1    g279(.A(G29gat), .ZN(new_n481));
  INV_X1    g280(.A(G36gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G50gat), .ZN(new_n487));
  INV_X1    g286(.A(G50gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G43gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n488), .B2(G43gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(KEYINPUT93), .A3(G50gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n501), .A3(new_n483), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n490), .B1(new_n502), .B2(new_n491), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n479), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n497), .A2(new_n493), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(new_n490), .A3(new_n491), .A4(new_n485), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(KEYINPUT17), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G15gat), .B(G22gat), .Z(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT95), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n510), .A2(KEYINPUT94), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT16), .B1(new_n514), .B2(G1gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G8gat), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n511), .A2(new_n519), .A3(new_n516), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n504), .A2(new_n508), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n511), .A2(new_n519), .A3(new_n516), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n519), .B1(new_n511), .B2(new_n516), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n523), .A2(new_n524), .B1(new_n498), .B2(new_n503), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n518), .A2(new_n505), .A3(new_n507), .A4(new_n520), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n525), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n522), .B(KEYINPUT13), .Z(new_n530));
  AOI21_X1  g329(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  AOI211_X1 g331(.A(KEYINPUT96), .B(new_n532), .C1(new_n528), .C2(new_n525), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n526), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n478), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n532), .B1(new_n528), .B2(new_n525), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n527), .ZN(new_n541));
  INV_X1    g340(.A(new_n478), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n537), .A4(new_n526), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT101), .ZN(new_n548));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  OR2_X1    g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(G85gat), .A3(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI221_X4 g360(.A(KEYINPUT102), .B1(new_n552), .B2(new_n553), .C1(new_n558), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT102), .ZN(new_n563));
  INV_X1    g362(.A(new_n552), .ZN(new_n564));
  NOR2_X1   g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n553), .A2(KEYINPUT102), .A3(new_n552), .ZN(new_n567));
  AND4_X1   g366(.A1(new_n566), .A2(new_n567), .A3(new_n558), .A4(new_n561), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n562), .A2(new_n568), .A3(KEYINPUT103), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n558), .A3(new_n561), .ZN(new_n570));
  INV_X1    g369(.A(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(new_n567), .A3(new_n558), .A4(new_n561), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT103), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n569), .A2(new_n504), .A3(new_n508), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT104), .ZN(new_n577));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n505), .A2(new_n507), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n580), .A2(new_n574), .B1(KEYINPUT41), .B2(new_n546), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n579), .B1(new_n577), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n551), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n578), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n550), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G57gat), .ZN(new_n590));
  INV_X1    g389(.A(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G57gat), .A2(G64gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT9), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  OR2_X1    g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  AND2_X1   g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n592), .A2(KEYINPUT97), .A3(new_n593), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n595), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT9), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n595), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n595), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n597), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n518), .B(new_n520), .C1(new_n611), .C2(new_n610), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT99), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT100), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n616), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n589), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n605), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n603), .A3(new_n602), .A4(new_n601), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n597), .B(new_n628), .C1(new_n562), .C2(new_n568), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n610), .A2(new_n572), .A3(new_n573), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(KEYINPUT105), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n610), .A2(new_n572), .A3(new_n634), .A4(new_n573), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n636), .B2(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n633), .B2(new_n635), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT106), .B1(new_n641), .B2(new_n631), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n633), .A2(new_n644), .A3(new_n635), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n645), .B1(new_n637), .B2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(new_n648), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n625), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n473), .A2(new_n544), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n465), .A2(new_n453), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n510), .ZN(G1324gat));
  OAI21_X1  g457(.A(G8gat), .B1(new_n655), .B2(new_n452), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n655), .A2(new_n452), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT107), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  AOI22_X1  g464(.A1(new_n663), .A2(new_n664), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667));
  AND4_X1   g466(.A1(new_n667), .A2(new_n662), .A3(new_n664), .A4(new_n665), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n666), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n305), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n655), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n459), .A2(G15gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n655), .B2(new_n672), .ZN(G1326gat));
  INV_X1    g472(.A(new_n426), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(G1327gat));
  NOR3_X1   g476(.A1(new_n589), .A2(new_n653), .A3(new_n624), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT109), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n473), .A2(new_n544), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n656), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n589), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n471), .A2(new_n472), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n456), .A2(KEYINPUT110), .A3(new_n426), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT110), .B1(new_n456), .B2(new_n426), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n691), .B2(new_n451), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n466), .B2(new_n674), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n451), .A2(new_n687), .A3(new_n694), .A4(new_n688), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n468), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n589), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n686), .B1(new_n699), .B2(new_n684), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n539), .A2(new_n543), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n653), .A2(new_n701), .A3(new_n624), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n656), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n703), .B2(new_n452), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n452), .A2(G36gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT46), .B1(new_n680), .B2(new_n708), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n680), .A2(KEYINPUT46), .A3(new_n708), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  OAI21_X1  g510(.A(new_n486), .B1(new_n680), .B2(new_n459), .ZN(new_n712));
  INV_X1    g511(.A(new_n468), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n451), .A2(new_n694), .A3(new_n688), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT111), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n715), .B2(new_n695), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n684), .B1(new_n716), .B2(new_n589), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n471), .A2(new_n472), .A3(new_n685), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n670), .A2(new_n486), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n702), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g521(.A1(new_n680), .A2(G50gat), .A3(new_n674), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n717), .A2(new_n426), .A3(new_n718), .A4(new_n702), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n723), .B2(new_n725), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(G1331gat));
  INV_X1    g528(.A(new_n653), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n625), .A2(new_n730), .A3(new_n544), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n697), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n656), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n590), .ZN(G1332gat));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n697), .A2(new_n731), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n445), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT49), .B(G64gat), .Z(new_n738));
  NOR3_X1   g537(.A1(new_n732), .A2(new_n452), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1333gat));
  NOR3_X1   g541(.A1(new_n732), .A2(G71gat), .A3(new_n459), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n305), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(G71gat), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n736), .A2(new_n426), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n715), .A2(new_n695), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n589), .B1(new_n750), .B2(new_n468), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n544), .A2(new_n624), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(new_n752), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n716), .A2(new_n754), .A3(new_n589), .A4(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n656), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n757), .A2(new_n559), .A3(new_n758), .A4(new_n653), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n730), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n700), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n656), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1336gat));
  NOR2_X1   g562(.A1(new_n452), .A2(G92gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n653), .B(new_n764), .C1(new_n753), .C2(new_n756), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n717), .A2(new_n445), .A3(new_n718), .A4(new_n760), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1337gat));
  NOR2_X1   g571(.A1(new_n459), .A2(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n653), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G99gat), .B1(new_n761), .B2(new_n670), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1338gat));
  NOR2_X1   g575(.A1(new_n674), .A2(G106gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n653), .B(new_n777), .C1(new_n753), .C2(new_n756), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n717), .A2(new_n426), .A3(new_n718), .A4(new_n760), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT53), .ZN(new_n782));
  INV_X1    g581(.A(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n779), .B2(KEYINPUT114), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n700), .A2(new_n785), .A3(new_n426), .A4(new_n760), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n787), .B2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(new_n624), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n640), .C1(new_n641), .C2(new_n631), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n651), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n794), .B2(new_n651), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n636), .A2(new_n630), .ZN(new_n799));
  INV_X1    g598(.A(new_n631), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n644), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n644), .B1(new_n803), .B2(KEYINPUT106), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n639), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n792), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n793), .B1(new_n637), .B2(new_n644), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n643), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(KEYINPUT55), .C1(new_n796), .C2(new_n797), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n806), .A2(new_n544), .A3(new_n649), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n522), .B1(new_n521), .B2(new_n525), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n529), .A2(new_n530), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n477), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n543), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n652), .B2(new_n649), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n698), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n649), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n585), .A2(new_n588), .A3(new_n543), .A4(new_n813), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n794), .A2(new_n651), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n795), .A3(new_n651), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n821), .A2(new_n822), .B1(new_n643), .B2(new_n807), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(KEYINPUT55), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n791), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n625), .A2(new_n544), .A3(new_n653), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n656), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n452), .A3(new_n460), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n701), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(new_n207), .ZN(G1340gat));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n730), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(new_n211), .ZN(G1341gat));
  NOR2_X1   g638(.A1(new_n835), .A2(new_n791), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(new_n218), .ZN(G1342gat));
  NOR2_X1   g640(.A1(new_n835), .A2(new_n589), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(KEYINPUT56), .A3(new_n227), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n842), .B2(new_n227), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n835), .B2(new_n589), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n305), .A2(new_n445), .A3(new_n674), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n834), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n544), .A2(new_n315), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n305), .A2(new_n656), .A3(new_n445), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n831), .B1(new_n826), .B2(new_n828), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n426), .ZN(new_n857));
  INV_X1    g656(.A(new_n819), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n643), .A2(new_n645), .A3(new_n648), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n823), .B2(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n860), .A3(new_n806), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n808), .B1(new_n796), .B2(new_n797), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n701), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n815), .B1(new_n864), .B2(new_n860), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(new_n698), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n791), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n674), .B1(new_n867), .B2(new_n828), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(new_n863), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n544), .B1(new_n823), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n816), .B1(new_n818), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n589), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n624), .B1(new_n874), .B2(new_n861), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n426), .C1(new_n875), .C2(new_n827), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT118), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n853), .B1(new_n857), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n701), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT58), .B1(new_n852), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n850), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(KEYINPUT58), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n853), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n869), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n827), .B1(new_n866), .B2(new_n791), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n889), .A4(new_n674), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n830), .A2(new_n426), .A3(new_n832), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n889), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT119), .B(new_n886), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n854), .A2(new_n855), .A3(new_n674), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n877), .B(new_n870), .C1(new_n896), .C2(KEYINPUT57), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n853), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G141gat), .B1(new_n900), .B2(new_n701), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n881), .B1(new_n885), .B2(new_n901), .ZN(G1344gat));
  NOR3_X1   g701(.A1(new_n848), .A2(G148gat), .A3(new_n730), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(KEYINPUT59), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n899), .B2(new_n653), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n426), .B1(new_n875), .B2(new_n827), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT122), .B1(new_n911), .B2(new_n889), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n892), .B2(new_n889), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n913), .A3(new_n653), .A4(new_n853), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n909), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT123), .B(new_n904), .C1(new_n908), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n879), .A2(KEYINPUT119), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n897), .A2(new_n895), .A3(new_n853), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n653), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n920), .B2(new_n906), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n921), .B2(new_n903), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n916), .A2(new_n922), .ZN(G1345gat));
  NOR2_X1   g722(.A1(new_n848), .A2(new_n791), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  AOI21_X1  g724(.A(G155gat), .B1(new_n924), .B2(KEYINPUT124), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n624), .A2(G155gat), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n925), .A2(new_n926), .B1(new_n899), .B2(new_n927), .ZN(G1346gat));
  INV_X1    g727(.A(new_n848), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n319), .B1(new_n929), .B2(new_n698), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n698), .A2(new_n319), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n899), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n833), .A2(new_n758), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n445), .A3(new_n460), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(G169gat), .A3(new_n701), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT125), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n656), .A2(new_n445), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(new_n459), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  OR3_X1    g738(.A1(new_n939), .A2(new_n426), .A3(new_n833), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n701), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n940), .B2(new_n730), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n653), .A2(new_n255), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n934), .B2(new_n944), .ZN(G1349gat));
  NOR3_X1   g744(.A1(new_n934), .A2(new_n268), .A3(new_n791), .ZN(new_n946));
  OR4_X1    g745(.A1(new_n426), .A2(new_n939), .A3(new_n791), .A4(new_n833), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G183gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n948), .B(new_n949), .ZN(G1350gat));
  OR2_X1    g749(.A1(new_n940), .A2(new_n589), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(G190gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n951), .B2(G190gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n698), .A2(new_n270), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n953), .A2(new_n954), .B1(new_n934), .B2(new_n955), .ZN(G1351gat));
  AND2_X1   g755(.A1(new_n910), .A2(new_n913), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n937), .A2(new_n305), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(G197gat), .A3(new_n544), .ZN(new_n960));
  INV_X1    g759(.A(G197gat), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n933), .A2(new_n445), .A3(new_n426), .A4(new_n670), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n701), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n960), .A2(new_n963), .ZN(G1352gat));
  NOR3_X1   g763(.A1(new_n962), .A2(G204gat), .A3(new_n730), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n957), .A2(new_n653), .A3(new_n958), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G204gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1353gat));
  OR3_X1    g768(.A1(new_n962), .A2(G211gat), .A3(new_n791), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n959), .A2(new_n624), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n698), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G218gat), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n589), .A2(G218gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n962), .B2(new_n977), .ZN(G1355gat));
endmodule


