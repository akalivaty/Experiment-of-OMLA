//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n208));
  OAI21_X1  g007(.A(G162gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218));
  AND4_X1   g017(.A1(new_n212), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n217), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n221), .A2(new_n215), .A3(new_n218), .A4(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n210), .A2(new_n219), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n231), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n224), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n220), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n216), .ZN(new_n246));
  NAND2_X1  g045(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n248), .B2(G162gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(G155gat), .B(G162gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n215), .A3(new_n218), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n243), .B(new_n240), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G141gat), .B(G148gat), .Z(new_n255));
  AOI21_X1  g054(.A(new_n211), .B1(new_n246), .B2(new_n247), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n250), .B(new_n255), .C1(new_n256), .C2(new_n244), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(KEYINPUT74), .A3(new_n240), .A4(new_n243), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n232), .A2(new_n236), .A3(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(new_n227), .C1(new_n230), .C2(new_n231), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n260), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n242), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G228gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT74), .B1(new_n224), .B2(new_n240), .ZN(new_n272));
  AND4_X1   g071(.A1(KEYINPUT74), .A2(new_n257), .A3(new_n240), .A4(new_n243), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n238), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n260), .A2(new_n263), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n238), .A3(new_n263), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n240), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n243), .B1(new_n249), .B2(new_n251), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n271), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n267), .A2(new_n271), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G22gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n206), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n266), .B2(new_n259), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n241), .B1(new_n274), .B2(new_n278), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n287), .B(new_n285), .C1(new_n288), .C2(new_n270), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n284), .B2(new_n285), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n270), .B1(new_n279), .B2(new_n242), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n270), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n254), .A2(new_n258), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n299), .A2(new_n238), .B1(new_n276), .B2(new_n277), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT81), .B(G22gat), .C1(new_n296), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n267), .A2(new_n271), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n303), .A2(KEYINPUT80), .A3(new_n285), .A4(new_n287), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n293), .A2(new_n295), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n291), .B1(new_n305), .B2(new_n205), .ZN(new_n306));
  INV_X1    g105(.A(G134gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G127gat), .ZN(new_n308));
  INV_X1    g107(.A(G127gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G113gat), .ZN(new_n315));
  INV_X1    g114(.A(G113gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT26), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(new_n326), .B2(KEYINPUT26), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  OR2_X1    g131(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(KEYINPUT28), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n332), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT27), .B(G183gat), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT67), .A4(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n336), .A3(G183gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT27), .B1(new_n338), .B2(KEYINPUT66), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n331), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n355), .A2(G169gat), .A3(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n326), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n323), .A2(KEYINPUT24), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n338), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(KEYINPUT23), .B2(new_n329), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(new_n356), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n333), .A2(new_n334), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n362), .B1(new_n372), .B2(G183gat), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n366), .A2(new_n367), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n322), .B1(new_n354), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT25), .A3(new_n358), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n326), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(KEYINPUT23), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n359), .A2(new_n361), .B1(new_n338), .B2(new_n363), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n313), .A2(new_n321), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n341), .A2(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n331), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT68), .ZN(new_n392));
  XOR2_X1   g191(.A(G71gat), .B(G99gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n387), .B1(new_n375), .B2(new_n385), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(KEYINPUT33), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n387), .A3(new_n385), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT34), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n375), .A2(new_n385), .A3(new_n399), .A4(new_n387), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n394), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n389), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n400), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n390), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  INV_X1    g207(.A(new_n390), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n306), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT71), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n382), .B1(new_n384), .B2(new_n331), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n238), .ZN(new_n422));
  INV_X1    g221(.A(new_n354), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(new_n382), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n422), .A2(new_n424), .A3(new_n266), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n238), .B1(new_n354), .B2(new_n374), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n419), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n420), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n278), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n418), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n266), .B1(new_n422), .B2(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n278), .A3(new_n428), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n417), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(KEYINPUT30), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n418), .C1(new_n425), .C2(new_n429), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n383), .B1(KEYINPUT3), .B2(new_n282), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n299), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n299), .A2(KEYINPUT75), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n282), .A2(new_n322), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(KEYINPUT4), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT77), .B1(new_n282), .B2(new_n322), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n224), .A2(new_n383), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(KEYINPUT4), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT76), .Z(new_n452));
  XOR2_X1   g251(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n443), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n446), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n444), .B2(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n441), .B2(new_n442), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT79), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n446), .B(new_n448), .C1(new_n224), .C2(new_n383), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n452), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n454), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n458), .A2(new_n459), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n299), .A2(KEYINPUT75), .A3(new_n438), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT75), .B1(new_n299), .B2(new_n438), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n453), .B1(new_n463), .B2(new_n452), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT79), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n456), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT0), .ZN(new_n475));
  XNOR2_X1  g274(.A(G57gat), .B(G85gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n477), .A2(KEYINPUT6), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n473), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n462), .B1(new_n461), .B2(new_n465), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT79), .A3(new_n471), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(new_n479), .A3(new_n456), .A4(new_n478), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n437), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n202), .B1(new_n413), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n407), .A2(new_n202), .A3(new_n411), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n306), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT82), .B1(new_n492), .B2(new_n489), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n489), .A3(KEYINPUT82), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n434), .A2(new_n436), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n480), .B(new_n482), .C1(new_n487), .C2(new_n456), .ZN(new_n497));
  INV_X1    g296(.A(new_n488), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n306), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  INV_X1    g300(.A(new_n411), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n407), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n450), .B1(new_n468), .B2(new_n469), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n452), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n463), .A2(new_n452), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT39), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n478), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n510), .A3(new_n452), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n512), .A2(KEYINPUT40), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT40), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n496), .B1(new_n473), .B2(new_n478), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n306), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT37), .B1(new_n425), .B2(new_n429), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT37), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n431), .A2(new_n520), .A3(new_n432), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n418), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT38), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT38), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n430), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n484), .A3(new_n488), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n506), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n494), .A2(new_n495), .B1(new_n500), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT13), .Z(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  AND2_X1   g332(.A1(KEYINPUT83), .A2(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT16), .B1(KEYINPUT83), .B2(G1gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(G1gat), .B2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI221_X1 g339(.A(new_n536), .B1(new_n537), .B2(new_n532), .C1(G1gat), .C2(new_n533), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  INV_X1    g346(.A(G36gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(KEYINPUT14), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(new_n546), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n553), .C1(new_n547), .C2(new_n548), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT15), .A3(new_n544), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n541), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n557), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT87), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT86), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n566), .A3(new_n561), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n531), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n558), .A2(KEYINPUT17), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n542), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n579), .A2(new_n580), .B1(G229gat), .B2(G233gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(new_n564), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n564), .A3(new_n581), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n569), .A2(new_n574), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n559), .A2(new_n562), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(new_n565), .A3(new_n567), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n590), .A2(new_n531), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT88), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n574), .A4(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n583), .ZN(new_n595));
  INV_X1    g394(.A(new_n574), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n529), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n601), .A2(KEYINPUT97), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT95), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n558), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  AOI211_X1 g414(.A(new_n602), .B(new_n614), .C1(KEYINPUT41), .C2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n575), .A3(new_n577), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n601), .A2(KEYINPUT97), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n616), .B(new_n619), .C1(KEYINPUT97), .C2(new_n601), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n624), .B(new_n627), .Z(new_n628));
  OR2_X1    g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT91), .B(G57gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G64gat), .ZN(new_n636));
  INV_X1    g435(.A(G64gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(G57gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n637), .A2(G57gat), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT89), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n629), .A2(new_n643), .A3(new_n630), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n629), .B2(new_n630), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT90), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT90), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n642), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n639), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n560), .B1(new_n653), .B2(KEYINPUT21), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT94), .Z(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(KEYINPUT21), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT92), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n659), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n639), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n604), .A2(new_n609), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT98), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n647), .A2(KEYINPUT90), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n651), .B1(new_n650), .B2(new_n642), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n669), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n612), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n612), .A3(new_n671), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT10), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n653), .A2(KEYINPUT10), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n613), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n668), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n668), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n676), .A2(new_n682), .A3(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n683), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n628), .A2(new_n667), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n600), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n497), .A2(new_n498), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g498(.A1(new_n695), .A2(new_n496), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n532), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n704), .B(new_n705), .C1(new_n532), .C2(new_n700), .ZN(G1325gat));
  NOR3_X1   g505(.A1(new_n695), .A2(G15gat), .A3(new_n412), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n696), .A2(new_n506), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(G15gat), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT100), .ZN(G1326gat));
  INV_X1    g509(.A(new_n306), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n667), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n692), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n628), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n600), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n547), .A3(new_n697), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n529), .B2(new_n628), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n306), .A2(new_n412), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT35), .B1(new_n723), .B2(new_n499), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n492), .A2(new_n489), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT82), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n727), .A3(new_n495), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n528), .A2(new_n500), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n624), .B(new_n627), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(KEYINPUT44), .A3(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n597), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT101), .B1(new_n594), .B2(new_n597), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n716), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n697), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n720), .A2(new_n741), .ZN(G1328gat));
  OAI21_X1  g541(.A(G36gat), .B1(new_n739), .B2(new_n496), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n718), .A2(new_n548), .A3(new_n437), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n743), .B(new_n747), .C1(new_n745), .C2(new_n744), .ZN(G1329gat));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n506), .A3(new_n732), .A4(new_n738), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G43gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n412), .A2(G43gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n718), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n752), .A3(KEYINPUT47), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n750), .A2(KEYINPUT103), .B1(new_n718), .B2(new_n751), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n755), .A3(G43gat), .ZN(new_n756));
  AOI211_X1 g555(.A(KEYINPUT104), .B(KEYINPUT47), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(KEYINPUT103), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n756), .A3(new_n752), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n753), .B1(new_n757), .B2(new_n762), .ZN(G1330gat));
  NAND4_X1  g562(.A1(new_n722), .A2(new_n306), .A3(new_n732), .A4(new_n738), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n711), .A2(G50gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n730), .A2(new_n598), .A3(new_n717), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT106), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n764), .A2(G50gat), .B1(KEYINPUT105), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n766), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n768), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT107), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n774), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n777));
  INV_X1    g576(.A(new_n772), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n765), .A3(new_n769), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(G1331gat));
  NOR2_X1   g580(.A1(new_n736), .A2(new_n692), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n667), .A3(new_n628), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n529), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n697), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(new_n635), .Z(G1332gat));
  XNOR2_X1  g585(.A(new_n496), .B(KEYINPUT108), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT109), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1333gat));
  INV_X1    g592(.A(new_n784), .ZN(new_n794));
  INV_X1    g593(.A(new_n506), .ZN(new_n795));
  OAI21_X1  g594(.A(G71gat), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n412), .A2(G71gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n306), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g601(.A1(new_n730), .A2(new_n715), .A3(new_n731), .A4(new_n737), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT51), .Z(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(new_n607), .A3(new_n697), .A4(new_n691), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n782), .A2(new_n715), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n733), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G85gat), .B1(new_n808), .B2(new_n740), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(G1336gat));
  NAND3_X1  g609(.A1(new_n787), .A2(new_n608), .A3(new_n691), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT111), .Z(new_n812));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(new_n804), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT112), .B1(new_n808), .B2(new_n788), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G92gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n808), .A2(KEYINPUT112), .A3(new_n788), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  OAI21_X1  g617(.A(G92gat), .B1(new_n808), .B2(new_n496), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n812), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n818), .B2(new_n821), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n808), .B2(new_n795), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n692), .A2(new_n412), .A3(G99gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1338gat));
  NOR3_X1   g625(.A1(new_n711), .A2(new_n692), .A3(G106gat), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n722), .A2(new_n306), .A3(new_n732), .A4(new_n807), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n804), .A2(new_n827), .B1(G106gat), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n828), .B2(G106gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT53), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n829), .B(new_n831), .ZN(G1339gat));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT10), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n674), .A2(new_n675), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n612), .B1(new_n653), .B2(new_n671), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n680), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n682), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(new_n681), .A3(KEYINPUT54), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n688), .B1(new_n681), .B2(KEYINPUT54), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n682), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n687), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n681), .A3(KEYINPUT54), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n842), .A2(new_n690), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n734), .A2(new_n735), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n590), .A2(new_n531), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n530), .B1(new_n578), .B2(new_n564), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n573), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n594), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n691), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n735), .ZN(new_n856));
  INV_X1    g655(.A(new_n848), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n597), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n691), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n855), .A2(new_n628), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n731), .A2(new_n857), .A3(new_n853), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n667), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n693), .A2(new_n736), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n306), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n740), .A2(new_n412), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n788), .A3(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n316), .A3(new_n599), .ZN(new_n871));
  INV_X1    g670(.A(new_n870), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n736), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n873), .B2(new_n316), .ZN(G1340gat));
  AND2_X1   g673(.A1(KEYINPUT115), .A2(G120gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(KEYINPUT115), .A2(G120gat), .ZN(new_n876));
  OAI22_X1  g675(.A1(new_n870), .A2(new_n692), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n691), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n875), .ZN(G1341gat));
  NOR2_X1   g678(.A1(new_n870), .A2(new_n715), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(new_n309), .ZN(G1342gat));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n869), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n731), .A2(new_n307), .A3(new_n496), .ZN(new_n883));
  XOR2_X1   g682(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G134gat), .B1(new_n870), .B2(new_n628), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G1343gat));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n306), .C1(new_n865), .C2(new_n866), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n795), .A2(new_n697), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n787), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n861), .B1(new_n599), .B2(new_n848), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n628), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n667), .B1(new_n897), .B2(new_n864), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n306), .B1(new_n898), .B2(new_n866), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n890), .B1(new_n901), .B2(new_n599), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n892), .A2(new_n900), .A3(KEYINPUT120), .A4(new_n598), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(G141gat), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n306), .B1(new_n865), .B2(new_n866), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n598), .A2(new_n213), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT118), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n895), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n900), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n736), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n908), .B1(new_n915), .B2(G141gat), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(G1344gat));
  NOR2_X1   g717(.A1(new_n711), .A2(KEYINPUT57), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n898), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n694), .A2(new_n599), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n692), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(KEYINPUT121), .B2(new_n895), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n923), .B(new_n925), .C1(new_n905), .C2(KEYINPUT57), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT59), .B1(new_n926), .B2(new_n214), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n912), .A2(new_n691), .A3(new_n914), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n214), .A2(KEYINPUT59), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n905), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n931), .A2(new_n214), .A3(new_n691), .A4(new_n894), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1345gat));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n914), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n248), .B1(new_n934), .B2(new_n715), .ZN(new_n935));
  OR4_X1    g734(.A1(new_n248), .A2(new_n905), .A3(new_n715), .A4(new_n895), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1346gat));
  OAI21_X1  g736(.A(G162gat), .B1(new_n934), .B2(new_n628), .ZN(new_n938));
  NOR4_X1   g737(.A1(new_n893), .A2(new_n628), .A3(G162gat), .A4(new_n437), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1347gat));
  OR2_X1    g741(.A1(new_n865), .A2(new_n866), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n697), .A2(new_n496), .A3(new_n412), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n711), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(new_n324), .A3(new_n599), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n788), .A2(new_n723), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n740), .B(new_n947), .C1(new_n865), .C2(new_n866), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n736), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n946), .A2(new_n950), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n945), .B2(new_n692), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n325), .A3(new_n691), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n715), .A2(new_n340), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n948), .A2(KEYINPUT123), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n948), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G183gat), .B1(new_n945), .B2(new_n715), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT60), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n344), .A3(new_n731), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n868), .A2(new_n731), .A3(new_n944), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(G190gat), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n967), .B2(G190gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  INV_X1    g771(.A(G197gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n795), .A2(new_n306), .A3(new_n787), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT124), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n943), .A2(new_n740), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n976), .B2(new_n737), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n923), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n506), .A2(new_n697), .A3(new_n496), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n599), .A2(new_n973), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n977), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n977), .B(KEYINPUT125), .C1(new_n980), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1352gat));
  XOR2_X1   g786(.A(KEYINPUT126), .B(G204gat), .Z(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(new_n980), .B2(new_n692), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n692), .A2(new_n989), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(KEYINPUT62), .B1(new_n976), .B2(new_n992), .ZN(new_n993));
  OR3_X1    g792(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n992), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(G1353gat));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n667), .A3(new_n979), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OR2_X1    g797(.A1(new_n715), .A2(G211gat), .ZN(new_n999));
  OAI22_X1  g798(.A1(new_n997), .A2(new_n998), .B1(new_n976), .B2(new_n999), .ZN(G1354gat));
  INV_X1    g799(.A(G218gat), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n976), .A2(new_n628), .ZN(new_n1002));
  INV_X1    g801(.A(new_n980), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n731), .A2(G218gat), .ZN(new_n1004));
  XOR2_X1   g803(.A(new_n1004), .B(KEYINPUT127), .Z(new_n1005));
  AOI22_X1  g804(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(G1355gat));
endmodule


