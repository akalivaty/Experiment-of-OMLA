

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U548 ( .A(n722), .B(n721), .ZN(n734) );
  BUF_X2 U549 ( .A(n887), .Z(n513) );
  XOR2_X1 U550 ( .A(KEYINPUT17), .B(n521), .Z(n887) );
  NOR2_X2 U551 ( .A1(n790), .A2(n679), .ZN(n695) );
  BUF_X1 U552 ( .A(n562), .Z(n553) );
  XOR2_X1 U553 ( .A(KEYINPUT14), .B(n577), .Z(n514) );
  NOR2_X1 U554 ( .A1(n766), .A2(n756), .ZN(n515) );
  XOR2_X1 U555 ( .A(n802), .B(KEYINPUT89), .Z(n516) );
  OR2_X1 U556 ( .A1(n695), .A2(n683), .ZN(n517) );
  XOR2_X1 U557 ( .A(KEYINPUT29), .B(n707), .Z(n518) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n717) );
  INV_X1 U559 ( .A(KEYINPUT101), .ZN(n721) );
  NAND2_X1 U560 ( .A1(n803), .A2(n516), .ZN(n804) );
  NOR2_X1 U561 ( .A1(G543), .A2(n537), .ZN(n530) );
  OR2_X1 U562 ( .A1(n805), .A2(n804), .ZN(n823) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n641) );
  NOR2_X1 U564 ( .A1(G651), .A2(n634), .ZN(n650) );
  XNOR2_X1 U565 ( .A(n529), .B(KEYINPUT64), .ZN(G160) );
  INV_X1 U566 ( .A(G2105), .ZN(n522) );
  AND2_X1 U567 ( .A1(n522), .A2(G2104), .ZN(n562) );
  AND2_X1 U568 ( .A1(G101), .A2(n562), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n519), .B(KEYINPUT23), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n520), .B(KEYINPUT65), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NAND2_X1 U572 ( .A1(G137), .A2(n513), .ZN(n526) );
  NOR2_X2 U573 ( .A1(G2104), .A2(n522), .ZN(n883) );
  NAND2_X1 U574 ( .A1(G125), .A2(n883), .ZN(n524) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U576 ( .A1(G113), .A2(n884), .ZN(n523) );
  AND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U580 ( .A(G651), .ZN(n537) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n530), .Z(n642) );
  NAND2_X1 U582 ( .A1(n642), .A2(G63), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT78), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  NAND2_X1 U585 ( .A1(G51), .A2(n650), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT79), .B(KEYINPUT6), .Z(n534) );
  XNOR2_X1 U588 ( .A(n535), .B(n534), .ZN(n543) );
  NAND2_X1 U589 ( .A1(n641), .A2(G89), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT4), .ZN(n539) );
  NOR2_X1 U591 ( .A1(n634), .A2(n537), .ZN(n645) );
  NAND2_X1 U592 ( .A1(G76), .A2(n645), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n540), .B(KEYINPUT77), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n541), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U597 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(G90), .A2(n641), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G77), .A2(n645), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G64), .A2(n642), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n650), .A2(G52), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT68), .B(n550), .Z(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U609 ( .A1(G99), .A2(n553), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G111), .A2(n884), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n883), .A2(G123), .ZN(n556) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n556), .Z(n557) );
  NOR2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n513), .A2(G135), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n929) );
  XNOR2_X1 U617 ( .A(G2096), .B(n929), .ZN(n561) );
  OR2_X1 U618 ( .A1(G2100), .A2(n561), .ZN(G156) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  INV_X1 U620 ( .A(G132), .ZN(G219) );
  INV_X1 U621 ( .A(G82), .ZN(G220) );
  NAND2_X1 U622 ( .A1(G102), .A2(n562), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G138), .A2(n513), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G126), .A2(n883), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G114), .A2(n884), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G164) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT72), .ZN(n570) );
  XNOR2_X1 U631 ( .A(KEYINPUT10), .B(n570), .ZN(G223) );
  INV_X1 U632 ( .A(G223), .ZN(n825) );
  NAND2_X1 U633 ( .A1(n825), .A2(G567), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n641), .A2(G81), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G68), .A2(n645), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n642), .A2(G56), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n514), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n650), .A2(G43), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n969) );
  XOR2_X1 U645 ( .A(G860), .B(KEYINPUT74), .Z(n601) );
  NOR2_X1 U646 ( .A1(n969), .A2(n601), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT75), .ZN(G153) );
  XOR2_X1 U648 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G92), .A2(n641), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G79), .A2(n645), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G66), .A2(n642), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G54), .A2(n650), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT15), .B(n588), .Z(n973) );
  INV_X1 U658 ( .A(n973), .ZN(n604) );
  INV_X1 U659 ( .A(G868), .ZN(n661) );
  NAND2_X1 U660 ( .A1(n604), .A2(n661), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G65), .A2(n642), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G53), .A2(n650), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT70), .B(n593), .Z(n595) );
  NAND2_X1 U666 ( .A1(n641), .A2(G91), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G78), .A2(n645), .ZN(n596) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n596), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n978) );
  XNOR2_X1 U671 ( .A(n978), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U672 ( .A1(G286), .A2(G868), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G299), .A2(n661), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U675 ( .A1(G559), .A2(n601), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT80), .B(n602), .Z(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT16), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT81), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n969), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G868), .A2(n973), .ZN(n607) );
  NOR2_X1 U682 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G559), .A2(n973), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n969), .B(n610), .ZN(n659) );
  NOR2_X1 U686 ( .A1(n659), .A2(G860), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G80), .A2(n645), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT82), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n641), .A2(G93), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G67), .A2(n642), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G55), .A2(n650), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n662) );
  XOR2_X1 U695 ( .A(n618), .B(n662), .Z(G145) );
  NAND2_X1 U696 ( .A1(G75), .A2(n645), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G62), .A2(n642), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G88), .A2(n641), .ZN(n621) );
  XNOR2_X1 U700 ( .A(KEYINPUT85), .B(n621), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n650), .A2(G50), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(G303) );
  NAND2_X1 U704 ( .A1(G72), .A2(n645), .ZN(n626) );
  XOR2_X1 U705 ( .A(KEYINPUT66), .B(n626), .Z(n631) );
  NAND2_X1 U706 ( .A1(G60), .A2(n642), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G47), .A2(n650), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT67), .B(n629), .Z(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n641), .A2(G85), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G49), .A2(n650), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n642), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n638) );
  XOR2_X1 U718 ( .A(KEYINPUT83), .B(n638), .Z(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G86), .A2(n641), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G61), .A2(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n645), .A2(G73), .ZN(n646) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(KEYINPUT84), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G48), .A2(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(G303), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G290), .ZN(n656) );
  XOR2_X1 U731 ( .A(n662), .B(G288), .Z(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(G299), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n658) );
  XNOR2_X1 U734 ( .A(G305), .B(KEYINPUT86), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n658), .B(n657), .ZN(n898) );
  XNOR2_X1 U736 ( .A(n898), .B(n659), .ZN(n660) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n664) );
  NOR2_X1 U738 ( .A1(G868), .A2(n662), .ZN(n663) );
  NOR2_X1 U739 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT87), .ZN(n666) );
  XNOR2_X1 U742 ( .A(KEYINPUT20), .B(n666), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U749 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G96), .A2(n672), .ZN(n831) );
  NAND2_X1 U751 ( .A1(n831), .A2(G2106), .ZN(n676) );
  NAND2_X1 U752 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U753 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(G69), .A2(n674), .ZN(n830) );
  NAND2_X1 U755 ( .A1(n830), .A2(G567), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n833) );
  NAND2_X1 U757 ( .A1(G661), .A2(G483), .ZN(n677) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n677), .ZN(n678) );
  NOR2_X1 U759 ( .A1(n833), .A2(n678), .ZN(n829) );
  NAND2_X1 U760 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U761 ( .A1(G40), .A2(G160), .ZN(n790) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n789) );
  INV_X1 U763 ( .A(n789), .ZN(n679) );
  OR2_X1 U764 ( .A1(n695), .A2(G1961), .ZN(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT25), .B(G2078), .ZN(n948) );
  NAND2_X1 U766 ( .A1(n695), .A2(n948), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n714) );
  NAND2_X1 U768 ( .A1(n714), .A2(G171), .ZN(n708) );
  AND2_X1 U769 ( .A1(n695), .A2(G1996), .ZN(n682) );
  XNOR2_X1 U770 ( .A(n682), .B(KEYINPUT26), .ZN(n686) );
  INV_X1 U771 ( .A(G1341), .ZN(n683) );
  INV_X1 U772 ( .A(n969), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n517), .A2(n684), .ZN(n685) );
  NOR2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n692) );
  NAND2_X1 U775 ( .A1(n692), .A2(n973), .ZN(n690) );
  INV_X1 U776 ( .A(n695), .ZN(n723) );
  NOR2_X1 U777 ( .A1(G2067), .A2(n723), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n695), .A2(G1348), .ZN(n687) );
  NOR2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n691), .B(KEYINPUT100), .ZN(n694) );
  OR2_X1 U782 ( .A1(n692), .A2(n973), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n695), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U785 ( .A(KEYINPUT27), .B(n696), .ZN(n699) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n723), .ZN(n697) );
  XOR2_X1 U787 ( .A(KEYINPUT98), .B(n697), .Z(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n978), .A2(n702), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U791 ( .A1(n978), .A2(n702), .ZN(n704) );
  XNOR2_X1 U792 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n703) );
  XNOR2_X1 U793 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n518), .ZN(n720) );
  NAND2_X1 U796 ( .A1(G8), .A2(n723), .ZN(n766) );
  NOR2_X1 U797 ( .A1(n766), .A2(G1966), .ZN(n709) );
  XNOR2_X1 U798 ( .A(n709), .B(KEYINPUT97), .ZN(n739) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n723), .ZN(n735) );
  INV_X1 U800 ( .A(n735), .ZN(n710) );
  AND2_X1 U801 ( .A1(G8), .A2(n710), .ZN(n711) );
  AND2_X1 U802 ( .A1(n739), .A2(n711), .ZN(n712) );
  XOR2_X1 U803 ( .A(n712), .B(KEYINPUT30), .Z(n713) );
  NOR2_X1 U804 ( .A1(G168), .A2(n713), .ZN(n716) );
  NOR2_X1 U805 ( .A1(G171), .A2(n714), .ZN(n715) );
  NOR2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U809 ( .A1(n734), .A2(G286), .ZN(n728) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n766), .ZN(n725) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U815 ( .A(n729), .B(KEYINPUT102), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n730), .A2(G8), .ZN(n733) );
  XOR2_X1 U817 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n731) );
  XNOR2_X1 U818 ( .A(KEYINPUT32), .B(n731), .ZN(n732) );
  XNOR2_X1 U819 ( .A(n733), .B(n732), .ZN(n742) );
  INV_X1 U820 ( .A(n734), .ZN(n738) );
  NAND2_X1 U821 ( .A1(G8), .A2(n735), .ZN(n736) );
  XOR2_X1 U822 ( .A(KEYINPUT96), .B(n736), .Z(n737) );
  NOR2_X1 U823 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U825 ( .A1(n742), .A2(n741), .ZN(n754) );
  NOR2_X1 U826 ( .A1(G2090), .A2(G303), .ZN(n743) );
  NAND2_X1 U827 ( .A1(G8), .A2(n743), .ZN(n744) );
  NAND2_X1 U828 ( .A1(n754), .A2(n744), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n745), .A2(n766), .ZN(n763) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n746) );
  XOR2_X1 U832 ( .A(n746), .B(KEYINPUT105), .Z(n747) );
  NOR2_X1 U833 ( .A1(n970), .A2(n747), .ZN(n748) );
  XNOR2_X1 U834 ( .A(n748), .B(KEYINPUT106), .ZN(n752) );
  XOR2_X1 U835 ( .A(G1981), .B(G305), .Z(n966) );
  INV_X1 U836 ( .A(n966), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n970), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n749), .A2(n766), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n757) );
  NAND2_X1 U840 ( .A1(n757), .A2(KEYINPUT33), .ZN(n755) );
  AND2_X1 U841 ( .A1(n752), .A2(n755), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n761) );
  INV_X1 U843 ( .A(n755), .ZN(n759) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n971) );
  INV_X1 U845 ( .A(n971), .ZN(n756) );
  AND2_X1 U846 ( .A1(n515), .A2(n757), .ZN(n758) );
  OR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n768) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U851 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n805) );
  NAND2_X1 U854 ( .A1(G105), .A2(n553), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(KEYINPUT38), .ZN(n776) );
  NAND2_X1 U856 ( .A1(G141), .A2(n513), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G117), .A2(n884), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G129), .A2(n883), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT93), .B(n772), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U863 ( .A(KEYINPUT94), .B(n777), .ZN(n863) );
  NAND2_X1 U864 ( .A1(G1996), .A2(n863), .ZN(n787) );
  NAND2_X1 U865 ( .A1(G131), .A2(n513), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT92), .ZN(n785) );
  NAND2_X1 U867 ( .A1(G95), .A2(n553), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G107), .A2(n884), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G119), .A2(n883), .ZN(n781) );
  XNOR2_X1 U871 ( .A(KEYINPUT91), .B(n781), .ZN(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n864) );
  NAND2_X1 U874 ( .A1(G1991), .A2(n864), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(KEYINPUT95), .B(n788), .ZN(n934) );
  INV_X1 U877 ( .A(n934), .ZN(n791) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n817) );
  NAND2_X1 U879 ( .A1(n791), .A2(n817), .ZN(n808) );
  NAND2_X1 U880 ( .A1(n513), .A2(G140), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(KEYINPUT90), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G104), .A2(n553), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n795), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G128), .A2(n883), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G116), .A2(n884), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT35), .B(n798), .Z(n799) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n801), .Z(n880) );
  XOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .Z(n816) );
  AND2_X1 U892 ( .A1(n880), .A2(n816), .ZN(n936) );
  NAND2_X1 U893 ( .A1(n936), .A2(n817), .ZN(n806) );
  AND2_X1 U894 ( .A1(n808), .A2(n806), .ZN(n803) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U896 ( .A1(n817), .A2(n984), .ZN(n802) );
  INV_X1 U897 ( .A(n806), .ZN(n821) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n863), .ZN(n807) );
  XOR2_X1 U899 ( .A(KEYINPUT107), .B(n807), .Z(n924) );
  INV_X1 U900 ( .A(n808), .ZN(n811) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n864), .ZN(n932) );
  NOR2_X1 U903 ( .A1(n809), .A2(n932), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n924), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(KEYINPUT108), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n817), .ZN(n819) );
  NOR2_X1 U909 ( .A1(n880), .A2(n816), .ZN(n941) );
  NAND2_X1 U910 ( .A1(n817), .A2(n941), .ZN(n818) );
  AND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  OR2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U914 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n825), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT110), .B(n826), .Z(n827) );
  NAND2_X1 U918 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n832), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n833), .ZN(G319) );
  XNOR2_X1 U929 ( .A(G1981), .B(KEYINPUT41), .ZN(n843) );
  XOR2_X1 U930 ( .A(G1986), .B(G1971), .Z(n835) );
  XNOR2_X1 U931 ( .A(G1961), .B(G1966), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U933 ( .A(G1991), .B(G1976), .Z(n837) );
  XNOR2_X1 U934 ( .A(G1956), .B(G1996), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2474), .B(KEYINPUT116), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n844), .B(KEYINPUT42), .ZN(n854) );
  XOR2_X1 U942 ( .A(KEYINPUT113), .B(G2100), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2678), .B(KEYINPUT114), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(G2096), .B(G2090), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT43), .B(KEYINPUT115), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U952 ( .A1(G124), .A2(n883), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT117), .B(n855), .Z(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G100), .A2(n553), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U957 ( .A1(G136), .A2(n513), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G112), .A2(n884), .ZN(n859) );
  NAND2_X1 U959 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U961 ( .A(n863), .B(G160), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n867) );
  XNOR2_X1 U964 ( .A(G164), .B(KEYINPUT121), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n869), .B(n868), .Z(n882) );
  NAND2_X1 U967 ( .A1(n513), .A2(G139), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n870), .B(KEYINPUT118), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G103), .A2(n553), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n873), .B(KEYINPUT119), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G127), .A2(n883), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G115), .A2(n884), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n876), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT120), .ZN(n919) );
  XNOR2_X1 U978 ( .A(n880), .B(n919), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n896) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U983 ( .A1(G106), .A2(n553), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G142), .A2(n513), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n893), .B(n929), .ZN(n894) );
  XNOR2_X1 U989 ( .A(G162), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n969), .B(n898), .ZN(n900) );
  XNOR2_X1 U993 ( .A(G171), .B(n973), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U995 ( .A(G286), .B(n901), .Z(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2430), .B(G2451), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2446), .B(G2427), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n911) );
  XOR2_X1 U1000 ( .A(G2438), .B(G2435), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G2443), .B(KEYINPUT109), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n907), .B(G2454), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  INV_X1 U1017 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n921) );
  XNOR2_X1 U1019 ( .A(G2072), .B(n919), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1021 ( .A(KEYINPUT50), .B(n922), .Z(n928) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n925), .Z(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT123), .B(n926), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n939) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT122), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n942), .ZN(n943) );
  XOR2_X1 U1036 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n962) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n962), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n944), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n957) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1041 ( .A1(n945), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n952) );
  XOR2_X1 U1045 ( .A(n948), .B(G27), .Z(n950) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G2084), .B(KEYINPUT54), .Z(n958) );
  XNOR2_X1 U1053 ( .A(G34), .B(n958), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1056 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n965), .ZN(n1019) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1060 ( .A(G168), .B(G1966), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n968), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1063 ( .A(n969), .B(G1341), .ZN(n987) );
  INV_X1 U1064 ( .A(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G166), .B(G1971), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n973), .B(G1348), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1070 ( .A(n978), .B(G1956), .Z(n980) );
  XOR2_X1 U1071 ( .A(G171), .B(G1961), .Z(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n1017) );
  INV_X1 U1079 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1080 ( .A(G1961), .B(KEYINPUT126), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(G5), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1085 ( .A(G1986), .B(G24), .Z(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1010) );
  XNOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(n1000), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(G1956), .B(G20), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1008), .Z(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

