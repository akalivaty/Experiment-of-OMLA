//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT3), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT81), .A2(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT81), .A2(G107), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT82), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT80), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT80), .A2(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT81), .B(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT82), .A3(new_n189), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n194), .A2(new_n199), .A3(new_n201), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT83), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n192), .A2(new_n193), .B1(new_n202), .B2(G107), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n208), .A2(new_n205), .A3(new_n201), .A4(new_n199), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n211), .B2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n217), .A3(new_n215), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT0), .B(G128), .Z(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n214), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n211), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n225), .A2(KEYINPUT0), .A3(G128), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n204), .A2(new_n231), .A3(new_n232), .A4(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n210), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n225), .A2(new_n235), .A3(G128), .A4(new_n227), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n226), .B1(new_n224), .B2(G146), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n241), .B(G101), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n242), .B2(new_n243), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT84), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n209), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n246), .A2(new_n244), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT10), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n226), .B2(new_n235), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n219), .A2(new_n221), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n209), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT11), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G134), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(G137), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n261), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n234), .A2(new_n249), .A3(new_n255), .A4(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT86), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n250), .A2(new_n209), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n236), .A3(new_n253), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n270), .B1(new_n280), .B2(new_n247), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n271), .A2(new_n283), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT87), .B(new_n276), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n234), .A2(new_n249), .A3(new_n255), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n257), .A2(new_n260), .B1(new_n256), .B2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n267), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n263), .B2(new_n289), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n284), .B2(new_n285), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n277), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n281), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n277), .B1(new_n302), .B2(new_n272), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n292), .B(new_n276), .C1(new_n284), .C2(new_n285), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(G469), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT9), .B(G234), .Z(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT74), .B(G125), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(KEYINPUT16), .A3(G140), .ZN(new_n314));
  INV_X1    g128(.A(new_n313), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(G125), .B2(G140), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n317), .B2(KEYINPUT16), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(G146), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n238), .A2(G119), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n238), .A2(G119), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G110), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n320), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n319), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n318), .A2(G146), .ZN(new_n330));
  XOR2_X1   g144(.A(G125), .B(G140), .Z(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n215), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n328), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n325), .B2(G110), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n333), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT22), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n329), .A2(new_n338), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(KEYINPUT77), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n297), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n312), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n346), .B2(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n312), .A3(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n297), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT79), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n343), .B2(new_n341), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n348), .A2(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n311), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n253), .A2(new_n236), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n256), .A2(KEYINPUT68), .A3(G137), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n256), .B2(G137), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT68), .B1(new_n256), .B2(G137), .ZN(new_n362));
  OAI21_X1  g176(.A(G131), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n290), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n291), .A2(new_n228), .A3(new_n223), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT2), .B(G113), .Z(new_n367));
  XNOR2_X1  g181(.A(G116), .B(G119), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT69), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n368), .B2(new_n367), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT28), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT67), .B1(new_n229), .B2(new_n270), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n291), .A2(new_n376), .A3(new_n228), .A4(new_n223), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n364), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n371), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(G101), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n274), .A3(G210), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n382), .B(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT30), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n371), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n372), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT31), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n385), .A4(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT71), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(KEYINPUT71), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n387), .B(new_n394), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(G472), .A2(G902), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n396), .B(KEYINPUT71), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n387), .A4(new_n394), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT32), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n401), .A2(new_n404), .A3(KEYINPUT32), .A4(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n405), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n391), .A2(new_n392), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n385), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n417), .C1(new_n380), .C2(new_n386), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n366), .A2(new_n371), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n374), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n385), .A2(KEYINPUT29), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n418), .B(new_n297), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G472), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n411), .A2(new_n413), .A3(new_n423), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n359), .A2(KEYINPUT89), .A3(new_n315), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT89), .B1(new_n359), .B2(new_n315), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n426), .C1(new_n230), .C2(new_n313), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n274), .A2(G224), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT90), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n427), .B(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(G110), .B(G122), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n371), .A2(new_n210), .A3(new_n233), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n369), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G113), .ZN(new_n436));
  INV_X1    g250(.A(G116), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n437), .A2(KEYINPUT5), .A3(G119), .ZN(new_n438));
  AOI211_X1 g252(.A(new_n436), .B(new_n438), .C1(KEYINPUT5), .C2(new_n368), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n250), .A3(new_n209), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n432), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n433), .A2(new_n441), .A3(new_n432), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n443), .A2(KEYINPUT88), .A3(KEYINPUT6), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n430), .B(new_n445), .C1(new_n446), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n428), .A2(KEYINPUT7), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n427), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n431), .B(KEYINPUT8), .Z(new_n453));
  INV_X1    g267(.A(new_n441), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n440), .B1(new_n209), .B2(new_n250), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n427), .A2(new_n451), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n452), .A2(new_n456), .A3(new_n457), .A4(new_n444), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n297), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n450), .A2(new_n297), .A3(new_n460), .A4(new_n458), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(KEYINPUT91), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n463), .A2(KEYINPUT91), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n468), .A2(G952), .A3(new_n274), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT21), .B(G898), .Z(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT97), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n319), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n383), .A2(new_n274), .A3(G214), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(G143), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n220), .A2(new_n478), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n264), .A4(new_n266), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n267), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n481), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT92), .B1(new_n488), .B2(KEYINPUT17), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(new_n483), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n477), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n188), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n333), .B1(new_n215), .B2(new_n317), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT18), .A2(G131), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n486), .A2(new_n495), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(KEYINPUT19), .B2(new_n317), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n330), .B(new_n488), .C1(new_n501), .C2(G146), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G475), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n297), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n499), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n493), .B1(new_n491), .B2(new_n498), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n297), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G475), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n507), .A4(new_n297), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n437), .A2(G122), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT95), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n437), .A2(G122), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n517), .B2(new_n518), .ZN(new_n523));
  OAI21_X1  g337(.A(G107), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n200), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT94), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n238), .A2(G143), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n220), .B2(new_n238), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G134), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n529), .A2(G134), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n524), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n308), .A2(new_n350), .A3(G953), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n530), .A2(KEYINPUT93), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n525), .B(new_n200), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT13), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n224), .A2(new_n536), .A3(G128), .ZN(new_n537));
  OAI211_X1 g351(.A(G134), .B(new_n537), .C1(new_n529), .C2(new_n536), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n530), .A2(KEYINPUT93), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n533), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n533), .B1(new_n532), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n297), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT96), .B(new_n297), .C1(new_n542), .C2(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n548), .B2(new_n544), .ZN(new_n551));
  NOR4_X1   g365(.A1(new_n467), .A2(new_n476), .A3(new_n516), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n358), .A2(new_n424), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT98), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  NAND3_X1  g369(.A1(new_n401), .A2(new_n297), .A3(new_n404), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G472), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n405), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n358), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n462), .A2(new_n463), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n465), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n476), .ZN(new_n563));
  INV_X1    g377(.A(new_n516), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n542), .A2(new_n543), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT33), .B1(new_n543), .B2(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n565), .A2(new_n566), .ZN(new_n569));
  OAI211_X1 g383(.A(G478), .B(new_n297), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n564), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n563), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n560), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n188), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n576), .B(new_n578), .ZN(G6));
  NAND4_X1  g393(.A1(new_n514), .A2(new_n510), .A3(new_n551), .A4(new_n515), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n562), .A2(new_n476), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n560), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G9));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n344), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n343), .B(new_n586), .Z(new_n587));
  AOI22_X1  g401(.A1(new_n348), .A2(new_n352), .B1(new_n354), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n552), .A2(new_n311), .A3(new_n559), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT37), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(G110), .Z(G12));
  OAI21_X1  g406(.A(new_n470), .B1(new_n472), .B2(G900), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n564), .A2(new_n551), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n562), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n589), .A2(new_n595), .A3(new_n309), .A4(new_n306), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n424), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G128), .ZN(G30));
  AOI21_X1  g413(.A(new_n412), .B1(new_n409), .B2(new_n410), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n414), .A2(new_n386), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n392), .A2(new_n419), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n386), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n604), .B2(new_n605), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT102), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n407), .A2(new_n408), .B1(KEYINPUT73), .B2(new_n405), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n611), .A2(new_n412), .A3(new_n612), .A4(new_n608), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n589), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n593), .B(KEYINPUT39), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n311), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(KEYINPUT40), .ZN(new_n618));
  INV_X1    g432(.A(new_n465), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n516), .A2(new_n551), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n464), .A2(new_n466), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT38), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(KEYINPUT40), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n615), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT103), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n220), .ZN(G45));
  AND3_X1   g441(.A1(new_n516), .A2(new_n572), .A3(new_n593), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n424), .A2(new_n597), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G146), .ZN(G48));
  INV_X1    g444(.A(new_n309), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n295), .A2(new_n297), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G469), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n298), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n287), .B2(new_n294), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(KEYINPUT104), .A3(new_n296), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n631), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n424), .A2(new_n575), .A3(new_n357), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT41), .B(G113), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G15));
  NAND4_X1  g455(.A1(new_n424), .A2(new_n357), .A3(new_n581), .A4(new_n638), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G116), .ZN(G18));
  NOR4_X1   g457(.A1(new_n588), .A2(new_n476), .A3(new_n516), .A4(new_n551), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n424), .A2(new_n595), .A3(new_n638), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G119), .ZN(G21));
  NAND2_X1  g460(.A1(new_n420), .A2(new_n386), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n403), .A2(new_n394), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n402), .B(KEYINPUT105), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n557), .A2(new_n357), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n557), .A2(new_n357), .A3(KEYINPUT106), .A4(new_n650), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n631), .B(new_n620), .C1(new_n634), .C2(new_n637), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n563), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G122), .ZN(G24));
  AND3_X1   g472(.A1(new_n589), .A2(new_n557), .A3(new_n650), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n638), .A3(new_n595), .A4(new_n628), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT107), .B(G125), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G27));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n303), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(KEYINPUT108), .B(new_n277), .C1(new_n302), .C2(new_n272), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(G469), .A3(new_n304), .A4(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT109), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT109), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n298), .A3(new_n300), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n309), .A2(new_n465), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n464), .B2(new_n466), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(KEYINPUT42), .A3(new_n628), .A4(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n407), .A2(new_n423), .A3(new_n408), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n357), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n669), .A2(new_n671), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n424), .A3(new_n357), .A4(new_n628), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n263), .ZN(G33));
  NAND4_X1  g494(.A1(new_n676), .A2(new_n424), .A3(new_n357), .A4(new_n594), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G134), .ZN(G36));
  NOR2_X1   g496(.A1(new_n516), .A2(new_n573), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(KEYINPUT43), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n686), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n685), .A2(KEYINPUT43), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n558), .A3(new_n589), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n664), .A2(KEYINPUT45), .A3(new_n304), .A4(new_n665), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n303), .A2(new_n304), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(G469), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT46), .B1(new_n699), .B2(new_n300), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(KEYINPUT46), .A3(new_n300), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n298), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n309), .A3(new_n616), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n692), .A2(new_n693), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n619), .B1(new_n464), .B2(new_n466), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G137), .ZN(G39));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n699), .A2(KEYINPUT46), .A3(new_n300), .ZN(new_n710));
  INV_X1    g524(.A(new_n298), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n700), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n709), .B1(new_n712), .B2(new_n631), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n703), .A2(KEYINPUT47), .A3(new_n309), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n628), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n357), .ZN(new_n717));
  INV_X1    g531(.A(new_n706), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n424), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G140), .ZN(G42));
  NAND4_X1  g535(.A1(new_n639), .A2(new_n642), .A3(new_n645), .A4(new_n657), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n516), .A2(new_n551), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n309), .A2(new_n589), .A3(new_n706), .A4(new_n306), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n424), .A2(new_n723), .A3(new_n593), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n676), .A2(new_n628), .A3(new_n659), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n681), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n580), .A2(KEYINPUT112), .B1(new_n516), .B2(new_n572), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n516), .A2(new_n572), .A3(KEYINPUT112), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n467), .A3(new_n476), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n358), .A2(new_n559), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n553), .A2(new_n732), .A3(new_n590), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n722), .A2(new_n679), .A3(new_n727), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n562), .A2(new_n620), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n309), .A2(new_n669), .A3(new_n588), .A4(new_n593), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n737), .C1(new_n610), .C2(new_n613), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n598), .A2(new_n629), .A3(new_n660), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n598), .A2(new_n629), .A3(new_n660), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT52), .A3(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n734), .A2(new_n744), .A3(KEYINPUT53), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT53), .B1(new_n734), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT54), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT113), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n298), .A2(KEYINPUT104), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n635), .A2(new_n296), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n309), .B(new_n595), .C1(new_n752), .C2(new_n636), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n589), .A2(new_n557), .A3(new_n628), .A4(new_n650), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n596), .B1(new_n600), .B2(new_n423), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n755), .B1(new_n594), .B2(new_n756), .ZN(new_n757));
  AND4_X1   g571(.A1(KEYINPUT52), .A2(new_n738), .A3(new_n757), .A4(new_n629), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(new_n742), .B2(new_n738), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n722), .A2(new_n733), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n679), .A2(new_n727), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n749), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n734), .A2(new_n744), .A3(KEYINPUT53), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT54), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n769), .A3(new_n765), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n764), .A2(KEYINPUT114), .A3(new_n769), .A4(new_n765), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n748), .A2(new_n768), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n715), .A2(KEYINPUT116), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n634), .A2(new_n637), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n631), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n713), .A2(new_n778), .A3(new_n714), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n470), .B1(new_n687), .B2(new_n690), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n655), .A2(new_n706), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n776), .A2(new_n671), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n469), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n614), .A2(new_n357), .A3(new_n789), .A4(new_n564), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n572), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n659), .A3(new_n781), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT117), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n623), .A2(new_n465), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n655), .A2(new_n638), .A3(new_n781), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n798), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(KEYINPUT50), .A3(new_n796), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n787), .A2(new_n794), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n712), .A2(new_n709), .A3(new_n631), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n703), .B2(new_n309), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n806), .B1(new_n809), .B2(new_n777), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n806), .A2(new_n713), .A3(new_n714), .A4(new_n777), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n810), .A2(new_n784), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n792), .B(KEYINPUT117), .Z(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n802), .C1(new_n572), .C2(new_n790), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n814), .B2(new_n803), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n805), .B1(new_n815), .B2(new_n786), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n798), .A2(new_n562), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT120), .ZN(new_n818));
  INV_X1    g632(.A(new_n674), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n788), .A2(new_n819), .A3(new_n781), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT48), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n614), .A2(new_n357), .A3(new_n789), .A4(new_n574), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(G952), .A3(new_n274), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n774), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n772), .A2(new_n773), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n767), .B1(new_n766), .B2(KEYINPUT54), .ZN(new_n828));
  AOI211_X1 g642(.A(KEYINPUT113), .B(new_n769), .C1(new_n764), .C2(new_n765), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n816), .A2(new_n818), .A3(new_n824), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n827), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(G952), .A2(G953), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n684), .A2(new_n670), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n836), .B(new_n357), .C1(new_n776), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n623), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n776), .A2(new_n837), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n614), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n835), .A2(new_n843), .ZN(G75));
  OAI211_X1 g658(.A(G210), .B(G902), .C1(new_n745), .C2(new_n746), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(KEYINPUT122), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT55), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n445), .B1(new_n446), .B2(new_n449), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n430), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(KEYINPUT122), .A3(new_n851), .A4(new_n846), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n848), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n274), .A2(G952), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G51));
  NAND2_X1  g670(.A1(new_n747), .A2(new_n770), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n300), .A2(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n300), .A2(KEYINPUT57), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(KEYINPUT123), .A3(new_n858), .A4(new_n859), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n295), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n766), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n297), .ZN(new_n866));
  INV_X1    g680(.A(new_n699), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n855), .B1(new_n864), .B2(new_n868), .ZN(G54));
  NAND3_X1  g683(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n870));
  INV_X1    g684(.A(new_n506), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n855), .ZN(G60));
  NOR2_X1   g688(.A1(new_n568), .A2(new_n569), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(G478), .A2(G902), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT59), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n774), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n857), .A2(new_n876), .A3(new_n878), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n855), .A3(new_n880), .ZN(G63));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n766), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n356), .B(KEYINPUT124), .Z(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n587), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n889), .A3(new_n855), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g705(.A1(new_n473), .A2(G224), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n761), .B2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n849), .B1(G898), .B2(new_n274), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(G69));
  NAND3_X1  g710(.A1(new_n704), .A2(new_n819), .A3(new_n736), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n681), .A2(new_n720), .A3(new_n707), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n679), .A2(new_n740), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n274), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n389), .A2(new_n390), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n501), .ZN(new_n902));
  INV_X1    g716(.A(G900), .ZN(new_n903));
  OAI21_X1  g717(.A(G953), .B1(new_n903), .B2(G227), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n626), .A2(new_n742), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n626), .A2(KEYINPUT62), .A3(new_n742), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n720), .A2(new_n707), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n424), .A2(new_n357), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n617), .A2(new_n912), .A3(new_n718), .A4(new_n730), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n274), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n902), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n915), .B2(new_n917), .ZN(G72));
  NAND3_X1  g732(.A1(new_n898), .A2(new_n761), .A3(new_n899), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n920));
  NAND2_X1  g734(.A1(G472), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n385), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n855), .B1(new_n924), .B2(new_n414), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT127), .Z(new_n926));
  INV_X1    g740(.A(new_n602), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n910), .A2(new_n761), .A3(new_n911), .A4(new_n913), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n923), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n922), .B(new_n865), .C1(new_n393), .C2(new_n416), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(G57));
endmodule


