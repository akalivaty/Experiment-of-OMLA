

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XOR2_X1 U324 ( .A(n377), .B(KEYINPUT18), .Z(n292) );
  AND2_X1 U325 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U326 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n376) );
  XOR2_X1 U327 ( .A(G120GAT), .B(G71GAT), .Z(n391) );
  XNOR2_X1 U328 ( .A(n322), .B(n293), .ZN(n323) );
  XNOR2_X1 U329 ( .A(n324), .B(n323), .ZN(n326) );
  NOR2_X1 U330 ( .A1(n546), .A2(n527), .ZN(n533) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n480) );
  XOR2_X1 U332 ( .A(n577), .B(KEYINPUT41), .Z(n551) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(n501) );
  XNOR2_X1 U334 ( .A(n480), .B(KEYINPUT58), .ZN(n481) );
  XNOR2_X1 U335 ( .A(n457), .B(G43GAT), .ZN(n458) );
  XNOR2_X1 U336 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n459), .B(n458), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n456) );
  XOR2_X1 U339 ( .A(G113GAT), .B(G36GAT), .Z(n295) );
  XNOR2_X1 U340 ( .A(G169GAT), .B(G50GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U342 ( .A(G8GAT), .B(G197GAT), .Z(n297) );
  XNOR2_X1 U343 ( .A(G141GAT), .B(G22GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n301) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT71), .B(n302), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U351 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n306) );
  XNOR2_X1 U352 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U354 ( .A(n308), .B(n307), .Z(n313) );
  XOR2_X1 U355 ( .A(G29GAT), .B(G43GAT), .Z(n310) );
  XNOR2_X1 U356 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n337) );
  XNOR2_X1 U358 ( .A(G15GAT), .B(G1GAT), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n311), .B(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U360 ( .A(n337), .B(n440), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n572) );
  INV_X1 U362 ( .A(G85GAT), .ZN(n314) );
  NAND2_X1 U363 ( .A1(G99GAT), .A2(n314), .ZN(n317) );
  INV_X1 U364 ( .A(G99GAT), .ZN(n315) );
  NAND2_X1 U365 ( .A1(n315), .A2(G85GAT), .ZN(n316) );
  NAND2_X1 U366 ( .A1(n317), .A2(n316), .ZN(n334) );
  XNOR2_X1 U367 ( .A(n391), .B(n334), .ZN(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U370 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n321) );
  XNOR2_X1 U371 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U373 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n325), .B(KEYINPUT13), .ZN(n439) );
  XOR2_X1 U375 ( .A(n326), .B(n439), .Z(n333) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n409) );
  XOR2_X1 U379 ( .A(G92GAT), .B(G64GAT), .Z(n330) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U382 ( .A(G204GAT), .B(n331), .Z(n379) );
  XNOR2_X1 U383 ( .A(n409), .B(n379), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n577) );
  NOR2_X1 U385 ( .A1(n572), .A2(n577), .ZN(n486) );
  XOR2_X1 U386 ( .A(G134GAT), .B(KEYINPUT80), .Z(n363) );
  XOR2_X1 U387 ( .A(n363), .B(n334), .Z(n336) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n416) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .Z(n385) );
  XNOR2_X1 U390 ( .A(n416), .B(n385), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U392 ( .A(G92GAT), .B(n337), .Z(n339) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(n341), .B(n340), .Z(n349) );
  XOR2_X1 U396 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n343) );
  XNOR2_X1 U397 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U399 ( .A(KEYINPUT79), .B(KEYINPUT65), .Z(n345) );
  XNOR2_X1 U400 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n557) );
  INV_X1 U404 ( .A(n557), .ZN(n479) );
  XOR2_X1 U405 ( .A(KEYINPUT36), .B(KEYINPUT105), .Z(n350) );
  XNOR2_X1 U406 ( .A(n479), .B(n350), .ZN(n585) );
  XOR2_X1 U407 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n352) );
  XNOR2_X1 U408 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(G141GAT), .B(n353), .Z(n420) );
  XOR2_X1 U411 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U414 ( .A(G57GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G1GAT), .B(G148GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n371) );
  XOR2_X1 U418 ( .A(G85GAT), .B(G162GAT), .Z(n361) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(G120GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U421 ( .A(n363), .B(n362), .Z(n365) );
  NAND2_X1 U422 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U424 ( .A(n366), .B(KEYINPUT5), .Z(n369) );
  XNOR2_X1 U425 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n367), .B(G127GAT), .ZN(n394) );
  XNOR2_X1 U427 ( .A(n394), .B(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n420), .B(n372), .ZN(n521) );
  INV_X1 U431 ( .A(n521), .ZN(n505) );
  XOR2_X1 U432 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n374) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U435 ( .A(n375), .B(KEYINPUT96), .Z(n381) );
  XNOR2_X1 U436 ( .A(n376), .B(KEYINPUT19), .ZN(n377) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(G183GAT), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n292), .B(n378), .ZN(n402) );
  XNOR2_X1 U439 ( .A(n402), .B(n379), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U441 ( .A(G8GAT), .B(KEYINPUT81), .Z(n444) );
  XOR2_X1 U442 ( .A(n382), .B(n444), .Z(n387) );
  XOR2_X1 U443 ( .A(G211GAT), .B(KEYINPUT21), .Z(n384) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(G218GAT), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n408) );
  XNOR2_X1 U446 ( .A(n408), .B(n385), .ZN(n386) );
  XNOR2_X2 U447 ( .A(n387), .B(n386), .ZN(n523) );
  XOR2_X1 U448 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n389) );
  XNOR2_X1 U449 ( .A(G134GAT), .B(G190GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U451 ( .A(n390), .B(G99GAT), .Z(n393) );
  XNOR2_X1 U452 ( .A(G43GAT), .B(n391), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U454 ( .A(n394), .B(G15GAT), .Z(n396) );
  NAND2_X1 U455 ( .A1(G227GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n404) );
  XOR2_X1 U458 ( .A(G176GAT), .B(KEYINPUT88), .Z(n400) );
  XNOR2_X1 U459 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n525) );
  NAND2_X1 U463 ( .A1(n523), .A2(n525), .ZN(n421) );
  XOR2_X1 U464 ( .A(KEYINPUT93), .B(KEYINPUT22), .Z(n406) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U467 ( .A(n407), .B(KEYINPUT92), .Z(n411) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U470 ( .A(G204GAT), .B(KEYINPUT89), .Z(n413) );
  XNOR2_X1 U471 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U473 ( .A(n415), .B(n414), .Z(n418) );
  XOR2_X1 U474 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XNOR2_X1 U475 ( .A(n416), .B(n443), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n476) );
  NAND2_X1 U478 ( .A1(n421), .A2(n476), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT101), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n423), .B(KEYINPUT25), .ZN(n427) );
  NOR2_X1 U481 ( .A1(n525), .A2(n476), .ZN(n425) );
  XNOR2_X1 U482 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n570) );
  XNOR2_X1 U484 ( .A(n523), .B(KEYINPUT27), .ZN(n429) );
  NAND2_X1 U485 ( .A1(n570), .A2(n429), .ZN(n426) );
  NAND2_X1 U486 ( .A1(n427), .A2(n426), .ZN(n428) );
  NAND2_X1 U487 ( .A1(n505), .A2(n428), .ZN(n432) );
  NAND2_X1 U488 ( .A1(n521), .A2(n429), .ZN(n546) );
  XOR2_X1 U489 ( .A(KEYINPUT28), .B(n476), .Z(n527) );
  XOR2_X1 U490 ( .A(n533), .B(KEYINPUT99), .Z(n430) );
  INV_X1 U491 ( .A(n525), .ZN(n535) );
  NAND2_X1 U492 ( .A1(n430), .A2(n535), .ZN(n431) );
  NAND2_X1 U493 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n433), .B(KEYINPUT102), .ZN(n484) );
  XOR2_X1 U495 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n435) );
  XNOR2_X1 U496 ( .A(G211GAT), .B(G64GAT), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n452) );
  XOR2_X1 U498 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n437) );
  NAND2_X1 U499 ( .A1(G231GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U501 ( .A(n438), .B(KEYINPUT15), .Z(n442) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n448) );
  XOR2_X1 U504 ( .A(n444), .B(n443), .Z(n446) );
  XNOR2_X1 U505 ( .A(G127GAT), .B(G71GAT), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U507 ( .A(n448), .B(n447), .Z(n450) );
  XNOR2_X1 U508 ( .A(G183GAT), .B(G78GAT), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U510 ( .A(n452), .B(n451), .Z(n581) );
  NAND2_X1 U511 ( .A1(n484), .A2(n581), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n585), .A2(n453), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT37), .B(n454), .Z(n518) );
  NAND2_X1 U514 ( .A1(n486), .A2(n518), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n501), .A2(n525), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n474) );
  XNOR2_X1 U518 ( .A(KEYINPUT64), .B(KEYINPUT116), .ZN(n472) );
  INV_X1 U519 ( .A(n572), .ZN(n547) );
  NAND2_X1 U520 ( .A1(n551), .A2(n547), .ZN(n461) );
  INV_X1 U521 ( .A(KEYINPUT46), .ZN(n460) );
  XOR2_X1 U522 ( .A(n461), .B(n460), .Z(n462) );
  NAND2_X1 U523 ( .A1(n462), .A2(n581), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n557), .A2(n463), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT47), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n585), .A2(n581), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT45), .B(n465), .Z(n466) );
  NOR2_X1 U528 ( .A1(n577), .A2(n466), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n467), .A2(n572), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n532) );
  NAND2_X1 U533 ( .A1(n532), .A2(n523), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n475), .A2(n521), .ZN(n571) );
  NAND2_X1 U536 ( .A1(n571), .A2(n476), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n525), .ZN(n567) );
  NOR2_X1 U539 ( .A1(n479), .A2(n567), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n557), .A2(n581), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n483), .ZN(n485) );
  AND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n504) );
  NAND2_X1 U544 ( .A1(n486), .A2(n504), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT103), .B(n487), .ZN(n494) );
  NAND2_X1 U546 ( .A1(n494), .A2(n521), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n494), .A2(n523), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U551 ( .A1(n494), .A2(n525), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n527), .A2(n494), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U556 ( .A1(n521), .A2(n501), .ZN(n498) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n523), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n527), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  INV_X1 U566 ( .A(n551), .ZN(n564) );
  NOR2_X1 U567 ( .A1(n547), .A2(n564), .ZN(n519) );
  NAND2_X1 U568 ( .A1(n519), .A2(n504), .ZN(n513) );
  NOR2_X1 U569 ( .A1(n505), .A2(n513), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  INV_X1 U573 ( .A(n523), .ZN(n509) );
  NOR2_X1 U574 ( .A1(n509), .A2(n513), .ZN(n510) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n535), .A2(n513), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(n511), .Z(n512) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  INV_X1 U579 ( .A(n527), .ZN(n514) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT114), .B(n520), .Z(n528) );
  NAND2_X1 U586 ( .A1(n521), .A2(n528), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .Z(n537) );
  NAND2_X1 U597 ( .A1(n532), .A2(n533), .ZN(n534) );
  NOR2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n547), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U602 ( .A1(n542), .A2(n551), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  INV_X1 U604 ( .A(n581), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n555), .A2(n542), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n557), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U612 ( .A1(n532), .A2(n570), .ZN(n545) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n558), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U618 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n558), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n572), .A2(n567), .ZN(n561) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n563) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n564), .A2(n567), .ZN(n565) );
  XOR2_X1 U632 ( .A(n566), .B(n565), .Z(G1349GAT) );
  NOR2_X1 U633 ( .A1(n581), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  XNOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n584) );
  NOR2_X1 U638 ( .A1(n572), .A2(n584), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n584), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

