//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT65), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n208), .B(new_n209), .C1(new_n205), .C2(new_n203), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n214), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n221));
  XOR2_X1   g020(.A(G183gat), .B(G190gat), .Z(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n203), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n220), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n225), .A2(new_n220), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n202), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n210), .A2(new_n218), .B1(new_n229), .B2(new_n235), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT69), .A3(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n237), .A2(new_n242), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT33), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n250));
  XOR2_X1   g049(.A(G15gat), .B(G43gat), .Z(new_n251));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n249), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n247), .B2(new_n248), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n247), .B2(new_n248), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n260), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n250), .B1(new_n249), .B2(new_n254), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n256), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n250), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n248), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(new_n269), .B2(new_n253), .ZN(new_n270));
  INV_X1    g069(.A(new_n263), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n270), .A2(new_n255), .B1(new_n271), .B2(new_n261), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n274), .B1(KEYINPUT22), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n237), .A2(KEYINPUT73), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n244), .B2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n244), .A2(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n244), .A2(KEYINPUT72), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n281), .B(new_n287), .C1(new_n290), .C2(new_n283), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n283), .A3(new_n289), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n237), .A2(new_n293), .A3(new_n282), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n294), .A3(new_n280), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n291), .A2(new_n295), .A3(new_n299), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(KEYINPUT30), .A3(new_n302), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n296), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT74), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G155gat), .B(G162gat), .Z(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n281), .B1(new_n315), .B2(new_n293), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n313), .B(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(G228gat), .B2(G233gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n311), .A2(new_n312), .ZN(new_n322));
  AOI211_X1 g121(.A(new_n321), .B(new_n316), .C1(new_n322), .C2(new_n318), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n320), .A2(G22gat), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(G22gat), .B1(new_n320), .B2(new_n323), .ZN(new_n326));
  XNOR2_X1  g125(.A(G78gat), .B(G106gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT31), .B(G50gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n326), .B1(new_n324), .B2(KEYINPUT79), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(G22gat), .C1(new_n320), .C2(new_n323), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n329), .B(KEYINPUT78), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n317), .A2(new_n242), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n241), .A2(new_n313), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT75), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n241), .B1(new_n313), .B2(new_n314), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n241), .B(new_n313), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n353), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n344), .B2(KEYINPUT4), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n343), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  INV_X1    g167(.A(new_n343), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n359), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT6), .B(new_n343), .C1(new_n360), .C2(new_n366), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT84), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(KEYINPUT35), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n273), .A2(new_n305), .A3(new_n338), .A4(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(KEYINPUT35), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n337), .B1(new_n265), .B2(new_n272), .ZN(new_n379));
  INV_X1    g178(.A(new_n377), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n305), .A3(new_n380), .A4(new_n375), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT80), .B(KEYINPUT39), .Z(new_n383));
  AND2_X1   g182(.A1(new_n355), .A2(new_n356), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n349), .B1(new_n344), .B2(new_n345), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n353), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n356), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n352), .B1(new_n351), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT39), .B1(new_n361), .B2(new_n353), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n386), .B(new_n369), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT40), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n390), .A2(KEYINPUT81), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n390), .B2(KEYINPUT81), .ZN(new_n393));
  INV_X1    g192(.A(new_n367), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n304), .A3(new_n303), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n395), .A2(new_n398), .A3(new_n304), .A4(new_n303), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n299), .B1(new_n291), .B2(new_n295), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT37), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n299), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n291), .B2(new_n295), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT38), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n372), .A2(new_n373), .A3(new_n302), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n280), .B(new_n287), .C1(new_n290), .C2(new_n283), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n292), .A2(new_n294), .A3(new_n281), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT37), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT38), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n296), .A2(KEYINPUT37), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n401), .B2(new_n403), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT83), .A3(KEYINPUT38), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n338), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n273), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n265), .A2(new_n272), .A3(KEYINPUT36), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n372), .A2(new_n373), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n338), .B1(new_n305), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n382), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G8gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(G1gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G1gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT16), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(new_n432), .A3(G8gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT14), .ZN(new_n441));
  INV_X1    g240(.A(G29gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n444));
  AOI21_X1  g243(.A(G36gat), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT15), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G36gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n444), .ZN(new_n450));
  NOR2_X1   g249(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT15), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n446), .ZN(new_n454));
  XNOR2_X1  g253(.A(G43gat), .B(G50gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(KEYINPUT15), .C1(new_n445), .C2(new_n447), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n456), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n440), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n437), .A2(new_n439), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT85), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT18), .ZN(new_n469));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(G197gat), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT11), .B(G169gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT12), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n464), .B(new_n465), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(new_n463), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n469), .A2(new_n474), .A3(new_n476), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT87), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n468), .A2(KEYINPUT18), .B1(new_n477), .B2(new_n479), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n474), .A4(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n476), .ZN(new_n487));
  INV_X1    g286(.A(new_n474), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n429), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G190gat), .B(G218gat), .Z(new_n493));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT41), .ZN(new_n495));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT8), .ZN(new_n499));
  NAND2_X1  g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G85gat), .ZN(new_n503));
  INV_X1    g302(.A(G92gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n499), .A2(new_n502), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n498), .ZN(new_n511));
  INV_X1    g310(.A(new_n498), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT92), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n512), .A2(new_n508), .ZN(new_n518));
  AOI22_X1  g317(.A1(KEYINPUT8), .A2(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n510), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n497), .B1(new_n465), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n460), .A2(new_n461), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n521), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n493), .A2(new_n494), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G134gat), .B(G162gat), .Z(new_n527));
  NAND2_X1  g326(.A1(new_n496), .A2(new_n495), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n526), .B(new_n529), .Z(new_n530));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  AND2_X1   g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G57gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G64gat), .ZN(new_n541));
  INV_X1    g340(.A(G64gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G57gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G78gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n538), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(new_n520), .A3(new_n514), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n517), .B2(new_n519), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n539), .B(new_n547), .C1(new_n552), .C2(new_n518), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n507), .A2(KEYINPUT94), .A3(new_n518), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n549), .B(new_n550), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n548), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n521), .A3(KEYINPUT10), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT95), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT97), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n560), .B1(new_n555), .B2(new_n557), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n533), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(KEYINPUT98), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n533), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT96), .B1(new_n572), .B2(new_n564), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n572), .A2(new_n564), .A3(KEYINPUT96), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n570), .A2(KEYINPUT98), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n548), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT20), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT89), .ZN(new_n587));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n583), .B(new_n584), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n464), .B1(KEYINPUT21), .B2(new_n556), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n590), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n590), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n578), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n593), .A3(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n577), .A3(new_n601), .ZN(new_n602));
  AOI211_X1 g401(.A(new_n530), .B(new_n576), .C1(new_n598), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n492), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n426), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n434), .ZN(G1324gat));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(new_n305), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT16), .B(G8gat), .Z(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(G8gat), .B1(new_n604), .B2(new_n305), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  MUX2_X1   g411(.A(new_n610), .B(new_n612), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g412(.A(G15gat), .B1(new_n607), .B2(new_n273), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n425), .A2(G15gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT99), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n607), .B2(new_n616), .ZN(G1326gat));
  XNOR2_X1  g416(.A(KEYINPUT43), .B(G22gat), .ZN(new_n618));
  OR3_X1    g417(.A1(new_n604), .A2(new_n338), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n604), .B2(new_n338), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(G1327gat));
  AND2_X1   g425(.A1(new_n397), .A2(new_n399), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n420), .A2(new_n338), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n428), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n382), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(KEYINPUT44), .A3(new_n530), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633));
  INV_X1    g432(.A(new_n530), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n429), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n426), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n598), .A2(new_n602), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n576), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n486), .A2(KEYINPUT102), .A3(new_n489), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT102), .B1(new_n486), .B2(new_n489), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n636), .A2(new_n637), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(G29gat), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n641), .A2(new_n634), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n492), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n442), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n652), .A2(new_n650), .A3(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(G1328gat));
  NOR2_X1   g455(.A1(new_n305), .A2(G36gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT46), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n652), .A2(KEYINPUT46), .A3(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n632), .A2(new_n635), .A3(new_n608), .A4(new_n647), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G36gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n659), .B(new_n660), .C1(new_n664), .C2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(new_n273), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n652), .A2(G43gat), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n632), .A2(new_n635), .A3(new_n425), .A4(new_n647), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G43gat), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n669), .B1(new_n668), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(G1330gat));
  NAND4_X1  g473(.A1(new_n632), .A2(new_n635), .A3(new_n337), .A4(new_n647), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G50gat), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT48), .B1(new_n676), .B2(KEYINPUT104), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n338), .A2(G50gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n492), .A2(new_n651), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n676), .B(new_n679), .C1(KEYINPUT104), .C2(KEYINPUT48), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1331gat));
  NOR4_X1   g482(.A1(new_n639), .A2(new_n645), .A3(new_n530), .A4(new_n640), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n631), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n426), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(new_n540), .ZN(G1332gat));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n305), .ZN(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  AND2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n688), .B2(new_n689), .ZN(G1333gat));
  INV_X1    g491(.A(G71gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n685), .B2(new_n667), .ZN(new_n694));
  INV_X1    g493(.A(new_n425), .ZN(new_n695));
  NOR4_X1   g494(.A1(new_n685), .A2(KEYINPUT105), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n631), .A2(new_n684), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n693), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n694), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g501(.A1(new_n698), .A2(new_n337), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g503(.A1(new_n426), .A2(G85gat), .A3(new_n640), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n638), .A2(new_n645), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n637), .B1(new_n304), .B2(new_n303), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n423), .B(new_n424), .C1(new_n707), .C2(new_n338), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT83), .B1(new_n418), .B2(KEYINPUT38), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n414), .B(new_n413), .C1(new_n401), .C2(new_n403), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n637), .A2(new_n710), .A3(new_n302), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n337), .B1(new_n712), .B2(new_n419), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n708), .B1(new_n713), .B2(new_n400), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n530), .B(new_n706), .C1(new_n714), .C2(new_n382), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n631), .A2(KEYINPUT51), .A3(new_n530), .A4(new_n706), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n705), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n576), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n636), .A2(new_n637), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n725), .B2(new_n503), .ZN(G1336gat));
  NAND4_X1  g525(.A1(new_n632), .A2(new_n635), .A3(new_n608), .A4(new_n724), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G92gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n305), .A2(new_n640), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n634), .B1(new_n629), .B2(new_n630), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT51), .B1(new_n730), .B2(new_n706), .ZN(new_n731));
  INV_X1    g530(.A(new_n706), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n429), .A2(new_n716), .A3(new_n634), .A4(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n504), .B(new_n729), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n728), .A2(new_n734), .A3(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT52), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n728), .A2(new_n734), .A3(KEYINPUT107), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1337gat));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n667), .A2(G99gat), .A3(new_n640), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT108), .Z(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT106), .B1(new_n731), .B2(new_n733), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n632), .A2(new_n635), .A3(new_n425), .A4(new_n724), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G99gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n740), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n720), .B2(new_n721), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1338gat));
  NAND4_X1  g552(.A1(new_n632), .A2(new_n635), .A3(new_n337), .A4(new_n724), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G106gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n338), .A2(G106gat), .A3(new_n640), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n731), .B2(new_n733), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n563), .A2(new_n760), .A3(new_n566), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n558), .B2(new_n561), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n555), .A2(new_n560), .A3(new_n557), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n533), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n574), .A2(new_n573), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(new_n764), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT111), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n774), .B(KEYINPUT55), .C1(new_n761), .C2(new_n764), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n768), .B(new_n770), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT112), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n490), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n564), .A2(new_n565), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT97), .B(new_n560), .C1(new_n555), .C2(new_n557), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n562), .A2(KEYINPUT54), .A3(new_n763), .ZN(new_n783));
  INV_X1    g582(.A(new_n533), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n772), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n774), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n771), .A2(KEYINPUT111), .A3(new_n772), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n789), .A2(new_n790), .A3(new_n770), .A4(new_n768), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n777), .A2(new_n779), .A3(new_n642), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n477), .A2(new_n479), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n473), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n486), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n640), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n530), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n486), .A2(new_n801), .A3(new_n795), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n530), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n777), .A2(new_n791), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n639), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n603), .A2(new_n646), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n337), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n305), .A2(new_n637), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n667), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n491), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT114), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n638), .A2(new_n634), .A3(new_n640), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n645), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n803), .A2(new_n804), .ZN(new_n817));
  INV_X1    g616(.A(new_n791), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n787), .A2(new_n788), .B1(new_n767), .B2(KEYINPUT110), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n790), .B1(new_n819), .B2(new_n770), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n797), .B1(new_n821), .B2(new_n645), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n817), .B1(new_n822), .B2(new_n530), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n816), .B1(new_n823), .B2(new_n639), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n426), .ZN(new_n825));
  INV_X1    g624(.A(new_n379), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n608), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(G113gat), .A3(new_n646), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n814), .A2(new_n829), .ZN(G1340gat));
  INV_X1    g629(.A(new_n828), .ZN(new_n831));
  AOI21_X1  g630(.A(G120gat), .B1(new_n831), .B2(new_n576), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n576), .A2(G120gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n811), .B2(new_n833), .ZN(G1341gat));
  NOR2_X1   g633(.A1(new_n828), .A2(new_n639), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n835), .B2(KEYINPUT115), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n638), .A2(G127gat), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n837), .B1(new_n811), .B2(new_n838), .ZN(G1342gat));
  OR3_X1    g638(.A1(new_n828), .A2(G134gat), .A3(new_n634), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n812), .B2(new_n634), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n846), .B(new_n847), .C1(new_n824), .C2(new_n338), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n338), .B1(new_n806), .B2(new_n807), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n849), .B2(KEYINPUT57), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n771), .B2(KEYINPUT117), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(KEYINPUT117), .B2(new_n771), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n490), .A2(new_n766), .A3(new_n765), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n634), .B1(new_n853), .B2(new_n797), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n638), .B1(new_n817), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT57), .B(new_n337), .C1(new_n855), .C2(new_n816), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n848), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n425), .A2(new_n809), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n645), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n425), .A2(new_n338), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n491), .A2(G141gat), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n825), .A2(new_n305), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n845), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n845), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n490), .A3(new_n858), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(G141gat), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT118), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(G141gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n865), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n825), .A2(new_n305), .A3(new_n861), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n859), .A2(G141gat), .B1(new_n873), .B2(new_n862), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n871), .B(new_n872), .C1(new_n874), .C2(new_n845), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n868), .A2(new_n875), .ZN(G1344gat));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n877), .A3(new_n576), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n849), .A2(KEYINPUT57), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n854), .B1(new_n776), .B2(new_n803), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n881), .A2(new_n639), .B1(new_n491), .B2(new_n603), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n847), .B1(new_n882), .B2(new_n338), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  MUX2_X1   g683(.A(new_n880), .B(new_n884), .S(KEYINPUT119), .Z(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n576), .A3(new_n858), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n857), .A2(new_n858), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n877), .C1(new_n888), .C2(new_n576), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n878), .B1(new_n887), .B2(new_n889), .ZN(G1345gat));
  INV_X1    g689(.A(G155gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n891), .A3(new_n638), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n888), .A2(new_n638), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n891), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n873), .B2(new_n530), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n530), .A2(G162gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(G1347gat));
  NAND2_X1  g696(.A1(new_n608), .A2(new_n426), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n667), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n808), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n491), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT121), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n824), .A2(new_n637), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n826), .A2(new_n305), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n646), .A2(G169gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  INV_X1    g709(.A(G176gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n901), .A2(new_n911), .A3(new_n640), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n908), .B2(new_n640), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n911), .C1(new_n908), .C2(new_n640), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n914), .B2(new_n916), .ZN(G1349gat));
  NAND4_X1  g716(.A1(new_n904), .A2(new_n211), .A3(new_n638), .A4(new_n905), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n808), .A2(new_n638), .A3(new_n899), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G183gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT125), .Z(new_n923));
  AOI21_X1  g722(.A(KEYINPUT123), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n919), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n921), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n925), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT124), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G1350gat));
  AOI21_X1  g728(.A(new_n212), .B1(new_n900), .B2(new_n530), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT61), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n530), .A2(new_n212), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n908), .B2(new_n932), .ZN(G1351gat));
  XOR2_X1   g732(.A(KEYINPUT126), .B(G197gat), .Z(new_n934));
  NOR2_X1   g733(.A1(new_n425), .A2(new_n898), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n885), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n936), .B2(new_n491), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n904), .A2(new_n861), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(new_n608), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n646), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(new_n941), .ZN(G1352gat));
  OAI21_X1  g741(.A(G204gat), .B1(new_n936), .B2(new_n640), .ZN(new_n943));
  INV_X1    g742(.A(G204gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n944), .A3(new_n729), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n939), .A2(new_n275), .A3(new_n638), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n885), .A2(new_n638), .A3(new_n935), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n936), .B2(new_n634), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n276), .A3(new_n530), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1355gat));
endmodule


