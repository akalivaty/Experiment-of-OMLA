//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n208), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT72), .B(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT71), .B(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n210), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT29), .B1(new_n208), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n230), .B2(new_n208), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n225), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n205), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n224), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n213), .A2(KEYINPUT29), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT78), .Z(new_n241));
  OR2_X1    g040(.A1(new_n229), .A2(new_n205), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n236), .B(new_n237), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n243), .A2(G22gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n204), .B1(new_n244), .B2(KEYINPUT79), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n243), .B(G22gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  OAI221_X1 g050(.A(new_n250), .B1(G183gat), .B2(G190gat), .C1(new_n251), .C2(KEYINPUT66), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(KEYINPUT66), .B2(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT23), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n258), .B2(new_n255), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n253), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n259), .A2(new_n261), .B1(new_n262), .B2(new_n251), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n261), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n266), .B2(new_n265), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT27), .B(G183gat), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT28), .Z(new_n272));
  AND2_X1   g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(G169gat), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(KEYINPUT26), .A3(new_n255), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n273), .B(new_n277), .C1(KEYINPUT26), .C2(new_n255), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G226gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n213), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n283), .B(new_n214), .C1(new_n280), .C2(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n291), .A3(new_n287), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n288), .A2(KEYINPUT30), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n299), .B2(new_n300), .ZN(new_n302));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n238), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT74), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n227), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n305), .A2(new_n306), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n308), .B2(KEYINPUT73), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n238), .B(new_n304), .ZN(new_n320));
  INV_X1    g119(.A(new_n312), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n309), .A2(new_n315), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n312), .B1(new_n309), .B2(new_n311), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT39), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT39), .B1(new_n320), .B2(new_n321), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n331), .B(new_n327), .C1(new_n329), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT40), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n334), .B2(new_n333), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n249), .B1(new_n298), .B2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n288), .A2(KEYINPUT37), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n291), .B1(new_n288), .B2(KEYINPUT37), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT38), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT38), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n327), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n344), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n328), .B2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n341), .A2(new_n294), .A3(new_n343), .A4(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n348), .A2(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(KEYINPUT76), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n328), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n328), .A2(new_n344), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n297), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n337), .A2(new_n350), .B1(new_n249), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n304), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n280), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n268), .A2(new_n360), .A3(new_n279), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT67), .A3(new_n364), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n363), .B2(KEYINPUT32), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n363), .B(KEYINPUT32), .C1(new_n364), .C2(new_n371), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n361), .A2(new_n359), .A3(new_n362), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT34), .B1(new_n359), .B2(KEYINPUT69), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n361), .A2(new_n362), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n358), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(KEYINPUT68), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n381), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n378), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n373), .B(new_n374), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT36), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n382), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n385), .A3(new_n374), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(KEYINPUT36), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n247), .A2(new_n248), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n383), .A2(new_n393), .A3(new_n387), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT35), .B1(new_n356), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n349), .A2(KEYINPUT35), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n297), .A4(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n357), .A2(new_n392), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G15gat), .ZN(new_n400));
  INV_X1    g199(.A(G15gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n402), .C1(new_n403), .C2(G1gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G22gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(G1gat), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G8gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT82), .B1(new_n405), .B2(G1gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI221_X1 g208(.A(new_n404), .B1(KEYINPUT82), .B2(G8gat), .C1(G1gat), .C2(new_n405), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g211(.A1(G29gat), .A2(G36gat), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(G43gat), .A2(G50gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(G43gat), .A2(G50gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(KEYINPUT15), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  NOR2_X1   g221(.A1(G43gat), .A2(G50gat), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT15), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(KEYINPUT80), .A2(G43gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(KEYINPUT80), .A2(G43gat), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n425), .A2(new_n426), .A3(G50gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT15), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n419), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n424), .B(new_n413), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n431));
  INV_X1    g230(.A(G36gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT81), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n415), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n412), .B(new_n421), .C1(new_n430), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR4_X1   g238(.A1(KEYINPUT81), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n414), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n420), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT80), .B(G43gat), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n428), .B(new_n419), .C1(new_n444), .C2(G50gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n412), .B1(new_n446), .B2(new_n421), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT83), .B(new_n411), .C1(new_n439), .C2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n409), .A2(new_n410), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n421), .B1(new_n430), .B2(new_n437), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT17), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n451), .B2(new_n438), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  INV_X1    g252(.A(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n411), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n448), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G229gat), .A2(G233gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT18), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n411), .B(new_n450), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n457), .B(KEYINPUT13), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n449), .A2(new_n450), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n454), .A2(new_n411), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT85), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n467), .A3(KEYINPUT84), .ZN(new_n468));
  XNOR2_X1  g267(.A(G113gat), .B(G141gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G197gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT11), .B(G169gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  XOR2_X1   g271(.A(new_n472), .B(KEYINPUT12), .Z(new_n473));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(new_n457), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n411), .B1(new_n439), .B2(new_n447), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT83), .B1(new_n449), .B2(new_n450), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(new_n448), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(KEYINPUT18), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n468), .B(new_n473), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n479), .A2(KEYINPUT18), .B1(new_n463), .B2(new_n466), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  INV_X1    g282(.A(new_n456), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n475), .ZN(new_n485));
  INV_X1    g284(.A(new_n473), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n482), .B(new_n485), .C1(KEYINPUT84), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n398), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(G71gat), .A2(G78gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G57gat), .B(G64gat), .Z(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(KEYINPUT9), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496));
  INV_X1    g295(.A(G57gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(G64gat), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n498), .A2(KEYINPUT87), .A3(G64gat), .A4(new_n499), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT88), .B1(new_n497), .B2(G64gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  INV_X1    g304(.A(G64gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(G57gat), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n492), .B1(new_n491), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n495), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT21), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n411), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G127gat), .B(G155gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT89), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n521), .A2(new_n523), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G183gat), .B(G211gat), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n521), .B(new_n523), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(new_n527), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n518), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n527), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n517), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G99gat), .B(G106gat), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n543), .A2(new_n544), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n549), .B2(new_n540), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n439), .B2(new_n447), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  AND2_X1   g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n450), .B1(KEYINPUT41), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT90), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n554), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n558), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n552), .A2(new_n564), .A3(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n564), .A4(new_n555), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n562), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(KEYINPUT92), .A3(new_n562), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n536), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n579));
  AND2_X1   g378(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT87), .B1(new_n582), .B2(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n511), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n495), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n553), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n512), .A2(new_n551), .A3(new_n586), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n553), .A2(KEYINPUT10), .A3(new_n512), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n578), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n578), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT94), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n577), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n490), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n355), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g407(.A(KEYINPUT16), .B(G8gat), .Z(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n298), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n610), .A2(KEYINPUT42), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(KEYINPUT42), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n298), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n613), .A2(KEYINPUT95), .A3(G8gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT95), .B1(new_n613), .B2(G8gat), .ZN(new_n615));
  OAI22_X1  g414(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(G1325gat));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n401), .A3(new_n391), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n392), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT96), .B(new_n388), .C1(new_n391), .C2(KEYINPUT36), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n605), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n622), .B2(new_n401), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(G1326gat));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n249), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT43), .B(G22gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  NOR3_X1   g427(.A1(new_n536), .A2(new_n576), .A3(new_n603), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n398), .A2(new_n489), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n632), .A2(G29gat), .A3(new_n355), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT45), .Z(new_n634));
  OAI21_X1  g433(.A(KEYINPUT44), .B1(new_n398), .B2(new_n576), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n357), .A2(new_n619), .A3(new_n620), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n395), .A2(new_n397), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n576), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT100), .B(new_n635), .C1(new_n640), .C2(KEYINPUT44), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n642), .B(KEYINPUT44), .C1(new_n398), .C2(new_n576), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n536), .B(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n481), .A2(KEYINPUT98), .A3(new_n487), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n481), .B2(new_n487), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n645), .A2(new_n603), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651), .B2(new_n355), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n652), .ZN(G1328gat));
  OAI21_X1  g452(.A(G36gat), .B1(new_n651), .B2(new_n297), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n631), .A2(new_n432), .A3(new_n298), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT46), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1329gat));
  NAND2_X1  g456(.A1(new_n621), .A2(new_n444), .ZN(new_n658));
  INV_X1    g457(.A(new_n391), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n632), .A2(new_n659), .ZN(new_n660));
  OAI22_X1  g459(.A1(new_n651), .A2(new_n658), .B1(new_n444), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g461(.A(G50gat), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n631), .A2(KEYINPUT101), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n249), .B1(new_n631), .B2(KEYINPUT101), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n393), .A2(new_n663), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n651), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g469(.A(new_n603), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n536), .A3(new_n576), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n671), .B(new_n672), .C1(new_n636), .C2(new_n637), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n606), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(new_n582), .Z(G1332gat));
  AOI21_X1  g474(.A(new_n297), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT102), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT103), .Z(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1333gat));
  NAND2_X1  g480(.A1(new_n673), .A2(new_n621), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n659), .A2(G71gat), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n682), .A2(G71gat), .B1(new_n673), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g484(.A1(new_n673), .A2(new_n249), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT104), .B(G78gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1335gat));
  NOR2_X1   g487(.A1(new_n648), .A2(new_n536), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n603), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n692));
  AOI211_X1 g491(.A(KEYINPUT44), .B(new_n576), .C1(new_n636), .C2(new_n637), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n643), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G85gat), .B1(new_n694), .B2(new_n355), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n638), .A2(new_n639), .A3(new_n689), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n671), .B1(new_n698), .B2(KEYINPUT105), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT105), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n606), .A2(new_n538), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(G1336gat));
  NOR3_X1   g501(.A1(new_n297), .A2(G92gat), .A3(new_n671), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT52), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n641), .A2(new_n298), .A3(new_n643), .A4(new_n691), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G92gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n703), .B(KEYINPUT106), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n705), .A2(G92gat), .B1(new_n698), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(G1337gat));
  XOR2_X1   g510(.A(KEYINPUT107), .B(G99gat), .Z(new_n712));
  INV_X1    g511(.A(new_n621), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n694), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n659), .A2(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n700), .B2(new_n715), .ZN(G1338gat));
  OAI21_X1  g515(.A(G106gat), .B1(new_n694), .B2(new_n393), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n393), .A2(G106gat), .A3(new_n671), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n717), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1339gat));
  NOR2_X1   g522(.A1(new_n672), .A2(new_n603), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n456), .A2(KEYINPUT110), .A3(new_n457), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT110), .B1(new_n456), .B2(new_n457), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n460), .A2(new_n462), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n472), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n603), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT10), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n587), .A2(new_n553), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n551), .B1(new_n512), .B2(new_n586), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n594), .A3(new_n591), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n593), .A3(KEYINPUT54), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n578), .B(new_n739), .C1(new_n590), .C2(new_n592), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n738), .A2(KEYINPUT55), .A3(new_n600), .A4(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n601), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n737), .A2(new_n593), .A3(KEYINPUT54), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n600), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n732), .B1(new_n649), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n576), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n730), .A2(new_n731), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n748), .A2(new_n576), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n725), .B1(new_n755), .B2(new_n645), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n355), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(new_n391), .A3(new_n393), .A4(new_n297), .ZN(new_n759));
  OAI21_X1  g558(.A(G113gat), .B1(new_n759), .B2(new_n489), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT112), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n757), .A2(new_n355), .A3(new_n298), .A4(new_n394), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n299), .A3(new_n648), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1340gat));
  NOR3_X1   g565(.A1(new_n759), .A2(new_n300), .A3(new_n671), .ZN(new_n767));
  AOI21_X1  g566(.A(G120gat), .B1(new_n762), .B2(new_n603), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1341gat));
  INV_X1    g568(.A(new_n645), .ZN(new_n770));
  OAI21_X1  g569(.A(G127gat), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(G127gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n772), .A3(new_n536), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1342gat));
  INV_X1    g573(.A(G134gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(new_n775), .A3(new_n639), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT56), .Z(new_n777));
  OAI21_X1  g576(.A(G134gat), .B1(new_n759), .B2(new_n576), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1343gat));
  NOR3_X1   g578(.A1(new_n621), .A2(new_n393), .A3(new_n298), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT116), .B1(new_n757), .B2(new_n355), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(G141gat), .A3(new_n489), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(KEYINPUT58), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n621), .A2(new_n355), .A3(new_n298), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788));
  INV_X1    g587(.A(new_n536), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n752), .A2(new_n754), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT114), .B1(new_n744), .B2(new_n745), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n738), .A2(new_n792), .A3(new_n600), .A4(new_n740), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n743), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n488), .A2(new_n794), .A3(new_n742), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n732), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n732), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n639), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n789), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n788), .B(new_n393), .C1(new_n801), .C2(new_n725), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n756), .B2(new_n249), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n787), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G141gat), .B1(new_n804), .B2(new_n489), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n804), .A2(new_n649), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n785), .B1(new_n808), .B2(G141gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(G1344gat));
  AOI21_X1  g609(.A(new_n788), .B1(new_n756), .B2(new_n249), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n249), .A2(new_n788), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n639), .A2(new_n813), .A3(new_n742), .A4(new_n746), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT118), .B1(new_n747), .B2(new_n576), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n750), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT119), .B1(new_n800), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n732), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT115), .B1(new_n795), .B2(new_n732), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n576), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(new_n816), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n789), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n577), .A2(new_n488), .A3(new_n603), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n812), .B1(new_n827), .B2(KEYINPUT120), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n811), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n603), .A3(new_n787), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(KEYINPUT121), .ZN(new_n833));
  OAI21_X1  g632(.A(G148gat), .B1(new_n832), .B2(KEYINPUT121), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT59), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(G148gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT59), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n804), .B2(new_n671), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n784), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n836), .A3(new_n603), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1345gat));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n215), .A3(new_n536), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n804), .A2(new_n770), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n215), .B2(new_n844), .ZN(G1346gat));
  OAI21_X1  g644(.A(G162gat), .B1(new_n804), .B2(new_n576), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n639), .A2(new_n216), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n784), .B2(new_n847), .ZN(G1347gat));
  NOR2_X1   g647(.A1(new_n606), .A2(new_n297), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n756), .A2(new_n391), .A3(new_n393), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G169gat), .B1(new_n850), .B2(new_n489), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n757), .A2(new_n606), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n394), .A2(new_n297), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n648), .A2(new_n274), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT122), .Z(G1348gat));
  OAI21_X1  g656(.A(G176gat), .B1(new_n850), .B2(new_n671), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n603), .A2(new_n275), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n854), .B2(new_n859), .ZN(G1349gat));
  INV_X1    g659(.A(new_n854), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n269), .A3(new_n536), .ZN(new_n862));
  OAI21_X1  g661(.A(G183gat), .B1(new_n850), .B2(new_n770), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n850), .B2(new_n576), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT61), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n270), .A3(new_n639), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1351gat));
  NAND3_X1  g668(.A1(new_n713), .A2(new_n249), .A3(new_n298), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n713), .A2(KEYINPUT123), .A3(new_n249), .A4(new_n298), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n649), .A2(G197gat), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n852), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n831), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n876), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n621), .A2(new_n606), .A3(new_n297), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n877), .A2(new_n488), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(G197gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT125), .B(new_n875), .C1(new_n880), .C2(G197gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(G1352gat));
  AND2_X1   g684(.A1(new_n873), .A2(new_n852), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n671), .A2(G204gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n872), .A3(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT62), .Z(new_n889));
  AND3_X1   g688(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n603), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G204gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(G1353gat));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n827), .A2(KEYINPUT120), .ZN(new_n895));
  INV_X1    g694(.A(new_n812), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n830), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n811), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n536), .A2(new_n619), .A3(new_n620), .A4(new_n849), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n897), .A2(KEYINPUT126), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G211gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT126), .B1(new_n831), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n900), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n886), .A2(new_n872), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n789), .A2(G211gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(KEYINPUT127), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1354gat));
  INV_X1    g715(.A(G218gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n909), .A2(new_n917), .A3(new_n639), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n890), .A2(new_n639), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(G1355gat));
endmodule


