//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT85), .ZN(new_n203));
  XOR2_X1   g002(.A(G78gat), .B(G106gat), .Z(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(KEYINPUT73), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n214), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n207), .A3(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n218), .B2(KEYINPUT73), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G141gat), .B(G148gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(G155gat), .B2(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G155gat), .B(G162gat), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT2), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n220), .B1(new_n238), .B2(KEYINPUT3), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n227), .A2(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n220), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G228gat), .ZN(new_n246));
  INV_X1    g045(.A(G233gat), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n241), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n240), .A2(KEYINPUT87), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n219), .B2(new_n239), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n219), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT86), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT86), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(new_n254), .C1(new_n219), .C2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n248), .B1(new_n253), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G22gat), .ZN(new_n263));
  INV_X1    g062(.A(G50gat), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n265), .B(new_n248), .C1(new_n253), .C2(new_n261), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n263), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n206), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G50gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n267), .A3(new_n205), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n242), .A2(new_n244), .ZN(new_n275));
  AND2_X1   g074(.A1(G113gat), .A2(G120gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(G113gat), .A2(G120gat), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT1), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT68), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n276), .B2(new_n277), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G113gat), .A2(G120gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n282), .A2(new_n287), .A3(new_n288), .A4(new_n279), .ZN(new_n289));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n288), .A3(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n294), .A3(new_n254), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n294), .A2(new_n238), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n242), .A2(new_n293), .A3(new_n289), .A4(new_n280), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n298), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT80), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n294), .A2(new_n238), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n296), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI211_X1 g110(.A(KEYINPUT80), .B(new_n296), .C1(new_n303), .C2(new_n308), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT5), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n314));
  NOR4_X1   g113(.A1(new_n294), .A2(new_n314), .A3(new_n238), .A4(KEYINPUT4), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n280), .A2(new_n289), .A3(new_n293), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n301), .B1(new_n316), .B2(new_n242), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n314), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n297), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n306), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G1gat), .B(G29gat), .Z(new_n322));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(KEYINPUT6), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n300), .A2(KEYINPUT79), .A3(new_n301), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n304), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT79), .B1(new_n300), .B2(new_n301), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n298), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(KEYINPUT5), .C1(new_n311), .C2(new_n312), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n326), .B1(new_n334), .B2(new_n306), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n326), .B(new_n306), .C1(new_n313), .C2(new_n320), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(KEYINPUT82), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(new_n340), .A3(new_n337), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n329), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G183gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT27), .B1(new_n343), .B2(KEYINPUT66), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(G183gat), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(G190gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n357));
  OAI22_X1  g156(.A1(new_n356), .A2(new_n357), .B1(new_n343), .B2(new_n348), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT67), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n348), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n345), .A2(G183gat), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n365), .B2(KEYINPUT27), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n366), .B2(new_n347), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n363), .B(new_n364), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT23), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(G183gat), .A3(G190gat), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n375), .A3(new_n377), .A4(new_n355), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n360), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n371), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n371), .B(KEYINPUT25), .C1(new_n378), .C2(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT74), .B1(new_n370), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n359), .A2(new_n369), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n219), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n383), .A2(new_n394), .A3(new_n384), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n395), .B2(new_n255), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n398), .B(new_n391), .C1(new_n395), .C2(new_n255), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n392), .B(new_n393), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n220), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n391), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n390), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n394), .A3(new_n391), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n219), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G8gat), .B(G36gat), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT77), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND3_X1  g208(.A1(new_n400), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n400), .A2(new_n412), .A3(new_n405), .A4(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n400), .A2(new_n405), .ZN(new_n415));
  INV_X1    g214(.A(new_n409), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT78), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n418), .B(new_n409), .C1(new_n400), .C2(new_n405), .ZN(new_n419));
  OAI22_X1  g218(.A1(new_n411), .A2(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n342), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n338), .A2(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n321), .A2(new_n327), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n341), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n328), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n415), .A2(new_n416), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n418), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n409), .B1(new_n400), .B2(new_n405), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n428), .A2(new_n430), .B1(new_n431), .B2(new_n413), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT83), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n274), .B1(new_n422), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n413), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(KEYINPUT88), .C1(new_n417), .C2(new_n419), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n296), .B1(new_n305), .B2(new_n295), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT39), .B1(new_n309), .B2(new_n310), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n327), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n424), .B1(new_n444), .B2(KEYINPUT40), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(KEYINPUT40), .B2(new_n444), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n274), .ZN(new_n448));
  INV_X1    g247(.A(new_n410), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n415), .A2(KEYINPUT37), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n416), .A2(KEYINPUT37), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n429), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n452), .B2(KEYINPUT38), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n335), .A2(new_n338), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n392), .B(new_n219), .C1(new_n397), .C2(new_n399), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n403), .A2(new_n393), .A3(new_n404), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(KEYINPUT37), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n463), .B(new_n464), .C1(new_n429), .C2(new_n451), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n429), .A2(new_n451), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT89), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n453), .A2(new_n457), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n448), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n316), .B1(new_n370), .B2(new_n385), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n387), .A2(new_n294), .A3(new_n388), .ZN(new_n471));
  INV_X1    g270(.A(G227gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n247), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n473), .B(KEYINPUT64), .Z(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  INV_X1    g278(.A(G15gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT32), .A3(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n477), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n471), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n472), .B2(new_n247), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n474), .A2(KEYINPUT34), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n490), .A2(KEYINPUT34), .B1(new_n492), .B2(KEYINPUT71), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n485), .A2(new_n493), .A3(new_n494), .A4(new_n487), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n496), .A2(new_n499), .A3(new_n497), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n434), .A2(new_n469), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n270), .A2(new_n273), .A3(new_n496), .A4(new_n497), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n421), .B1(new_n342), .B2(new_n420), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n426), .A2(new_n432), .A3(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n436), .B2(new_n438), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n507), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(G57gat), .A2(G64gat), .ZN(new_n519));
  AND2_X1   g318(.A1(G71gat), .A2(G78gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(KEYINPUT9), .ZN(new_n521));
  INV_X1    g320(.A(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT100), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n527), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(KEYINPUT21), .ZN(new_n531));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G127gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n541), .A2(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT94), .B(G8gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n543), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G8gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(KEYINPUT21), .B2(new_n530), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT101), .Z(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n234), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n553), .B(new_n555), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n557));
  OR3_X1    g356(.A1(new_n540), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n540), .B2(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT14), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(G29gat), .ZN(new_n573));
  INV_X1    g372(.A(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT14), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT91), .B(G36gat), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n572), .B(new_n575), .C1(new_n576), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n482), .A2(G50gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT15), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n264), .A2(G43gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n578), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT15), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n581), .A2(new_n583), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n570), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n568), .B(new_n569), .Z(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n592), .A2(new_n595), .B1(KEYINPUT102), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(KEYINPUT102), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  OR2_X1    g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT103), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n600), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n601), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n561), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n550), .A3(new_n548), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n551), .A2(new_n584), .A3(new_n586), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n551), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n591), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n589), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n620), .B(KEYINPUT96), .C1(new_n621), .C2(new_n589), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n613), .A3(new_n610), .A4(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT18), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G197gat), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT11), .B(G169gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n625), .A2(new_n610), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n613), .A4(new_n624), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n631), .A3(new_n618), .ZN(new_n641));
  INV_X1    g440(.A(new_n630), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n641), .B(new_n636), .C1(new_n642), .C2(new_n628), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n594), .A2(new_n528), .A3(new_n529), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n530), .A2(new_n570), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n647), .A2(new_n649), .A3(KEYINPUT104), .A4(new_n648), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n530), .A2(KEYINPUT10), .A3(new_n570), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n646), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n649), .ZN(new_n657));
  INV_X1    g456(.A(new_n646), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n656), .B2(new_n659), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n645), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(KEYINPUT105), .A3(new_n663), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n608), .A2(new_n644), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n517), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n342), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g473(.A1(new_n436), .A2(new_n438), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(G8gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT106), .Z(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n498), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n672), .A2(new_n480), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n672), .A2(new_n505), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n687), .B2(new_n480), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT107), .Z(G1326gat));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n274), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n607), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n644), .A2(new_n561), .A3(new_n670), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n517), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n573), .A3(new_n342), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n434), .A2(new_n469), .A3(new_n506), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n512), .A2(KEYINPUT35), .B1(new_n514), .B2(new_n515), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n517), .A2(KEYINPUT44), .A3(new_n693), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n694), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n426), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n697), .A2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n695), .A2(new_n676), .A3(new_n576), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n705), .A2(new_n675), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n576), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n505), .A2(G43gat), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n695), .A2(new_n685), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n705), .A2(new_n713), .B1(G43gat), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g515(.A1(new_n448), .A2(new_n264), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n703), .A3(new_n694), .A4(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n517), .A2(new_n274), .A3(new_n693), .A4(new_n694), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n264), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n718), .A2(KEYINPUT108), .A3(new_n719), .A4(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n718), .A2(new_n721), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT109), .B1(new_n727), .B2(KEYINPUT48), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n729), .B(new_n719), .C1(new_n718), .C2(new_n721), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n724), .A2(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n722), .A2(new_n723), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n725), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n734), .B(new_n735), .C1(new_n728), .C2(new_n730), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n638), .A2(new_n643), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n608), .A2(new_n738), .A3(new_n669), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n517), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n342), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743));
  INV_X1    g542(.A(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n676), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n744), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  NAND2_X1  g548(.A1(new_n740), .A2(new_n505), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n498), .A2(G71gat), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(G71gat), .B1(new_n740), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n274), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n561), .A2(new_n738), .A3(new_n669), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n704), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n426), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n700), .A2(new_n738), .A3(new_n561), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n761));
  OR2_X1    g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n670), .A2(new_n565), .A3(new_n342), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(G1336gat));
  INV_X1    g566(.A(new_n758), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n676), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G92gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n675), .A2(new_n669), .A3(G92gat), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(new_n764), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n760), .B(new_n774), .Z(new_n775));
  AOI22_X1  g574(.A1(new_n769), .A2(G92gat), .B1(new_n775), .B2(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n758), .B2(new_n506), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n670), .A2(new_n685), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n765), .B2(new_n781), .ZN(G1338gat));
  NAND2_X1  g581(.A1(new_n768), .A2(new_n274), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n448), .A2(new_n669), .A3(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n764), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n785), .B(KEYINPUT115), .Z(new_n788));
  AOI22_X1  g587(.A1(new_n783), .A2(G106gat), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(G1339gat));
  NAND4_X1  g590(.A1(new_n644), .A2(new_n561), .A3(new_n607), .A4(new_n669), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n653), .A2(new_n654), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n650), .A2(new_n651), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n658), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n656), .A2(new_n796), .A3(KEYINPUT54), .ZN(new_n797));
  INV_X1    g596(.A(new_n662), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n656), .B2(KEYINPUT54), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n793), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n658), .B1(new_n794), .B2(new_n795), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n662), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n656), .A2(new_n796), .A3(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n663), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n638), .B2(new_n643), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n630), .A2(new_n640), .A3(new_n618), .A4(new_n637), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n613), .B1(new_n639), .B2(new_n624), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n611), .A2(new_n615), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n635), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n808), .A2(new_n811), .A3(new_n668), .A4(new_n666), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n607), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n560), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n811), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n806), .B1(new_n815), .B2(KEYINPUT116), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n808), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n607), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n792), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n792), .B(new_n822), .C1(new_n814), .C2(new_n819), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n426), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n514), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n738), .A2(new_n283), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT118), .Z(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n823), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n342), .A3(new_n448), .A4(new_n675), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n498), .A3(new_n644), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n831), .B2(new_n283), .ZN(G1340gat));
  AOI21_X1  g631(.A(G120gat), .B1(new_n825), .B2(new_n670), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n830), .A2(new_n284), .A3(new_n780), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1341gat));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n534), .A3(new_n561), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n830), .A2(new_n498), .A3(new_n560), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n534), .ZN(G1342gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n607), .A2(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n514), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT119), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n842), .B2(KEYINPUT56), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n830), .A2(new_n498), .A3(new_n607), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n842), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1343gat));
  NOR3_X1   g650(.A1(new_n676), .A2(new_n505), .A3(new_n426), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n829), .B2(new_n274), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n820), .A2(new_n274), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n852), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G141gat), .B1(new_n859), .B2(new_n644), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n676), .A2(new_n505), .A3(new_n448), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n824), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n228), .A3(new_n738), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n860), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n230), .A3(new_n670), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT122), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n670), .B(new_n852), .C1(new_n855), .C2(new_n858), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n230), .A2(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(KEYINPUT123), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n816), .A2(new_n818), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n693), .ZN(new_n880));
  INV_X1    g679(.A(new_n806), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n738), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n607), .A2(new_n812), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n884), .A3(new_n560), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n822), .B1(new_n885), .B2(new_n792), .ZN(new_n886));
  INV_X1    g685(.A(new_n823), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n274), .B(new_n854), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n448), .B1(new_n821), .B2(new_n823), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT124), .A3(new_n854), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n856), .A2(new_n857), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n670), .A3(new_n852), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n878), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n870), .B1(new_n877), .B2(new_n896), .ZN(G1345gat));
  OAI21_X1  g696(.A(G155gat), .B1(new_n859), .B2(new_n560), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n862), .A2(new_n234), .A3(new_n561), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  NOR3_X1   g699(.A1(new_n859), .A2(new_n235), .A3(new_n607), .ZN(new_n901));
  AOI21_X1  g700(.A(G162gat), .B1(new_n862), .B2(new_n693), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n676), .A2(new_n426), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n821), .B2(new_n823), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n509), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n738), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(G169gat), .ZN(G1348gat));
  NAND4_X1  g707(.A1(new_n905), .A2(new_n448), .A3(new_n685), .A4(new_n670), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n561), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(new_n351), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n343), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1350gat));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n906), .A2(new_n693), .B1(new_n918), .B2(new_n348), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n348), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n505), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n891), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n738), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n922), .B(KEYINPUT126), .Z(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT127), .Z(new_n928));
  AND2_X1   g727(.A1(new_n894), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n738), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n923), .A2(G204gat), .A3(new_n669), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n894), .A2(new_n928), .A3(new_n670), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n925), .A2(new_n209), .A3(new_n561), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n927), .A2(new_n561), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n894), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  AOI211_X1 g740(.A(new_n941), .B(new_n209), .C1(new_n894), .C2(new_n938), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n937), .B1(new_n940), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n925), .B2(new_n693), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n607), .A2(new_n210), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n929), .B2(new_n945), .ZN(G1355gat));
endmodule


