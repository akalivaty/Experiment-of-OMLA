//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g049(.A(KEYINPUT66), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n469), .A3(G125), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n477), .A2(new_n469), .A3(KEYINPUT64), .A4(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  INV_X1    g061(.A(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n468), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n491), .A2(new_n468), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n493), .A2(KEYINPUT67), .A3(G124), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n493), .B2(G124), .ZN(new_n495));
  OAI221_X1 g070(.A(new_n488), .B1(new_n489), .B2(new_n490), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n477), .A3(new_n469), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT69), .B1(new_n468), .B2(G114), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(G126), .A2(G2105), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n491), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n498), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(G2105), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(KEYINPUT69), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(new_n508), .B1(new_n501), .B2(new_n502), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .ZN(new_n519));
  NAND2_X1  g094(.A1(G126), .A2(G2105), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n521), .A2(new_n465), .A3(new_n469), .A4(new_n467), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G164));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(G543), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n531), .A2(G651), .B1(new_n535), .B2(G50), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n532), .A2(new_n533), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n529), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT5), .B(G543), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n540), .B(KEYINPUT71), .C1(new_n533), .C2(new_n532), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G88), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(G303));
  INV_X1    g119(.A(G303), .ZN(G166));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT7), .Z(new_n547));
  NAND3_X1  g122(.A1(new_n540), .A2(G63), .A3(G651), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n547), .B(new_n549), .C1(G51), .C2(new_n535), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n539), .A2(new_n541), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G89), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  NAND2_X1  g129(.A1(new_n551), .A2(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n529), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n535), .B2(G52), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G43), .B2(new_n535), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n551), .A2(G81), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n566), .B(new_n567), .C1(new_n565), .C2(new_n564), .ZN(new_n568));
  INV_X1    g143(.A(G860), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n568), .A2(new_n569), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT73), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n529), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n551), .A2(G91), .B1(G651), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT74), .B1(new_n534), .B2(new_n580), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(KEYINPUT9), .A3(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(G299));
  NAND2_X1  g164(.A1(new_n551), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n535), .A2(G49), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n539), .A2(new_n541), .A3(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n535), .A2(G48), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OR2_X1    g174(.A1(KEYINPUT5), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(KEYINPUT5), .A2(G543), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT77), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n605), .A2(G73), .A3(G543), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G651), .C1(new_n602), .C2(new_n607), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n598), .A2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n551), .A2(G85), .ZN(new_n614));
  NAND2_X1  g189(.A1(G72), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G60), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n529), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(new_n535), .B2(G47), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n542), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(G79), .A2(G543), .ZN(new_n626));
  INV_X1    g201(.A(G66), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n529), .B2(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n628), .A2(G651), .B1(new_n535), .B2(G54), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n620), .B1(new_n631), .B2(G868), .ZN(G284));
  XNOR2_X1  g207(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g208(.A1(G286), .A2(G868), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT80), .Z(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n631), .B1(new_n639), .B2(G860), .ZN(G148));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n568), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n630), .A2(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(new_n641), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g220(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n487), .A2(G135), .ZN(new_n650));
  OR2_X1    g225(.A1(G99), .A2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n651), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n652));
  INV_X1    g227(.A(G123), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n652), .C1(new_n492), .C2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT82), .B(G2438), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n660), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  INV_X1    g250(.A(G14), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n682), .B2(new_n679), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(new_n693), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n694), .A2(new_n696), .A3(new_n700), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT88), .Z(new_n711));
  OR3_X1    g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  OAI21_X1  g293(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(G286), .A2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n719), .B(KEYINPUT98), .S(new_n721), .Z(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G19), .B(new_n568), .S(G16), .Z(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G1341), .ZN(new_n726));
  NOR2_X1   g301(.A1(G171), .A2(new_n720), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G5), .B2(new_n720), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT30), .B(G28), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n734), .C1(new_n654), .C2(new_n733), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n728), .B2(new_n729), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n725), .A2(G1341), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(G32), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(new_n742), .B1(G105), .B2(new_n462), .ZN(new_n743));
  INV_X1    g318(.A(G129), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n492), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G141), .B2(new_n487), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(new_n733), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n730), .A2(new_n736), .A3(new_n737), .A4(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n724), .A2(new_n726), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n720), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT100), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT23), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n636), .B2(new_n720), .ZN(new_n756));
  INV_X1    g331(.A(G1956), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n733), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n752), .B(new_n758), .C1(G2084), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G162), .A2(G29), .ZN(new_n765));
  OR2_X1    g340(.A1(G29), .A2(G35), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT29), .B(G2090), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n733), .A2(G27), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n733), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT99), .B(G2078), .Z(new_n774));
  XOR2_X1   g349(.A(new_n773), .B(new_n774), .Z(new_n775));
  INV_X1    g350(.A(G1348), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n631), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n733), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT91), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT28), .ZN(new_n783));
  INV_X1    g358(.A(G128), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n468), .A2(G116), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n492), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n487), .A2(G140), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(new_n733), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G1348), .B2(new_n778), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n770), .A2(new_n771), .A3(new_n780), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n764), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G33), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT92), .Z(new_n796));
  NAND3_X1  g371(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  NAND3_X1  g374(.A1(new_n477), .A2(new_n469), .A3(G127), .ZN(new_n800));
  NAND2_X1  g375(.A1(G115), .A2(G2104), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G139), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n802), .A2(new_n468), .B1(new_n803), .B2(new_n470), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n796), .B1(new_n806), .B2(new_n733), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  INV_X1    g383(.A(G2072), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT95), .Z(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n763), .A2(G2084), .B1(new_n748), .B2(new_n749), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT97), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n811), .A2(new_n818), .A3(new_n813), .A4(new_n814), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n794), .A2(new_n816), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n794), .A2(new_n816), .A3(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT101), .ZN(new_n822));
  OR2_X1    g397(.A1(G6), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G305), .B2(new_n720), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1981), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n720), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n720), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1971), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n720), .A2(G23), .ZN(new_n833));
  INV_X1    g408(.A(G288), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n720), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT33), .B(G1976), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n826), .A2(new_n831), .A3(new_n832), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n840));
  MUX2_X1   g415(.A(G24), .B(G290), .S(G16), .Z(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G1986), .Z(new_n842));
  NOR2_X1   g417(.A1(G25), .A2(G29), .ZN(new_n843));
  INV_X1    g418(.A(G119), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n468), .A2(G107), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n492), .A2(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n487), .A2(G131), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n843), .B1(new_n849), .B2(G29), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G1991), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n842), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n840), .A2(KEYINPUT90), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT90), .B1(new_n840), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n839), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT36), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n839), .B(new_n859), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n820), .A2(new_n822), .B1(new_n858), .B2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n822), .A2(new_n820), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(G150));
  NOR2_X1   g439(.A1(new_n630), .A2(new_n639), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n529), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n869), .A2(G651), .B1(new_n535), .B2(G55), .ZN(new_n870));
  INV_X1    g445(.A(G93), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n542), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n568), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n568), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n866), .B(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n569), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(G860), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT102), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(G145));
  INV_X1    g458(.A(new_n789), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n518), .A2(new_n522), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n789), .B1(new_n522), .B2(new_n518), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n746), .ZN(new_n889));
  INV_X1    g464(.A(new_n746), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n805), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n806), .A3(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n849), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(new_n647), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n647), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n487), .A2(G142), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT103), .Z(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(G118), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n493), .B2(G130), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n898), .A2(new_n901), .A3(new_n905), .A4(new_n897), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT104), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT104), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n895), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n485), .B(new_n654), .Z(new_n913));
  XNOR2_X1  g488(.A(G162), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n893), .A2(new_n909), .A3(new_n894), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n914), .B1(new_n912), .B2(new_n915), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g498(.A(G305), .B(G288), .Z(new_n924));
  XNOR2_X1  g499(.A(G290), .B(G166), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT42), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n875), .B(new_n643), .Z(new_n929));
  OAI21_X1  g504(.A(new_n630), .B1(new_n587), .B2(new_n588), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n585), .A2(new_n586), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n585), .A2(new_n586), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n631), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT105), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND3_X1  g510(.A1(G299), .A2(new_n935), .A3(new_n631), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n927), .A2(new_n928), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n927), .A2(new_n928), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(KEYINPUT41), .A3(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n930), .A2(new_n933), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n929), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n939), .B1(new_n938), .B2(new_n945), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n872), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(G868), .B2(new_n950), .ZN(G295));
  INV_X1    g526(.A(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n641), .B1(new_n952), .B2(new_n946), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n950), .A2(G868), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n949), .B(new_n956), .C1(G868), .C2(new_n950), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(G331));
  OAI21_X1  g533(.A(G171), .B1(G286), .B2(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g534(.A1(G286), .A2(KEYINPUT108), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n873), .A2(new_n874), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n873), .B2(new_n874), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n874), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n568), .A2(new_n872), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT108), .B(G286), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n959), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n873), .A2(new_n874), .A3(new_n960), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n940), .A3(new_n942), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n963), .A2(new_n936), .A3(new_n969), .A4(new_n934), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n926), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n917), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n971), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(new_n926), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n971), .A2(new_n975), .A3(new_n972), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n930), .A2(new_n933), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT41), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n961), .A2(new_n962), .A3(new_n959), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n967), .B1(new_n966), .B2(new_n968), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT41), .B1(new_n934), .B2(new_n936), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n937), .A2(new_n941), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n970), .A4(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n972), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n926), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n973), .A2(new_n917), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n994), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n981), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n980), .B2(new_n998), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1001), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g577(.A(KEYINPUT125), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT114), .B(G8), .Z(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n524), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n885), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1009));
  INV_X1    g584(.A(G40), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n483), .B2(G2105), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(new_n1011), .A3(new_n474), .A4(new_n475), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT115), .B(G2084), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1008), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n484), .A2(new_n474), .A3(G40), .A4(new_n475), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT45), .B1(new_n885), .B2(new_n1007), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n524), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1966), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1005), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G168), .A2(new_n1004), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT51), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1007), .B1(new_n511), .B2(new_n514), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n476), .A2(new_n1027), .A3(new_n1011), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1026), .B(G1384), .C1(new_n515), .C2(new_n523), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n723), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT70), .B1(new_n518), .B2(new_n522), .ZN(new_n1031));
  AND4_X1   g606(.A1(KEYINPUT70), .A2(new_n522), .A3(new_n503), .A4(new_n510), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1007), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1016), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1036), .A3(new_n1013), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1030), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1022), .B1(new_n1038), .B2(G8), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1024), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1022), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1038), .A2(KEYINPUT122), .A3(new_n1022), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1041), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1011), .A2(new_n474), .A3(new_n475), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n518), .B2(new_n522), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT45), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1384), .B1(new_n515), .B2(new_n523), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1050), .B(new_n1052), .C1(KEYINPUT45), .C2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1054), .B2(G2078), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n729), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT123), .A4(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(KEYINPUT53), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1018), .A2(new_n1059), .A3(new_n1019), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n609), .A2(new_n611), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n596), .A2(new_n597), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1068), .A2(new_n1069), .A3(G1981), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n598), .B2(new_n612), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1067), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1011), .A2(new_n1051), .A3(new_n474), .A4(new_n475), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1004), .ZN(new_n1076));
  OAI21_X1  g651(.A(G1981), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n598), .A2(new_n1071), .A3(new_n612), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n834), .A2(G1976), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1076), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1005), .B(new_n1074), .C1(G288), .C2(new_n1082), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT55), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n524), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1050), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2090), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1033), .B2(new_n1026), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1971), .B1(new_n1095), .B2(new_n1050), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1005), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1087), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1089), .ZN(new_n1099));
  INV_X1    g674(.A(G1971), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1052), .B1(new_n1053), .B2(KEYINPUT45), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT113), .B(new_n1100), .C1(new_n1101), .C2(new_n1016), .ZN(new_n1102));
  INV_X1    g677(.A(G2090), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1034), .A2(new_n1036), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT113), .B1(new_n1054), .B2(new_n1100), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(new_n1099), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1066), .A2(new_n1098), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1003), .B1(new_n1048), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1022), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1112), .A2(new_n1024), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1113), .A2(new_n1042), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1041), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1090), .A2(new_n1050), .A3(new_n1091), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1116), .A2(new_n1103), .B1(new_n1054), .B2(new_n1100), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1089), .B1(new_n1117), .B2(new_n1004), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1080), .A2(new_n1086), .A3(new_n1084), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1107), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n1120), .A3(KEYINPUT125), .A4(new_n1066), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1109), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G301), .B(KEYINPUT54), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1016), .A2(KEYINPUT124), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n1059), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1017), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1016), .A2(KEYINPUT124), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1058), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1057), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1123), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1113), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT56), .B(G2072), .Z(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n1054), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1135), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1095), .A2(new_n1137), .A3(new_n1050), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1092), .A2(new_n757), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n585), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n579), .A2(KEYINPUT57), .A3(new_n583), .A4(new_n584), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT61), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1136), .A2(KEYINPUT120), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1144), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n1153), .B2(new_n1145), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n776), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1155));
  INV_X1    g730(.A(G2067), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1075), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1155), .A2(new_n630), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n630), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT60), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1016), .A2(G1996), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  AOI22_X1  g737(.A1(new_n1095), .A2(new_n1161), .B1(new_n1074), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1164), .A2(KEYINPUT121), .ZN(new_n1165));
  OR3_X1    g740(.A1(new_n1163), .A2(new_n568), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n630), .A2(KEYINPUT60), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1155), .A2(new_n1167), .A3(new_n1157), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1164), .A2(KEYINPUT121), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1165), .B(new_n1169), .C1(new_n1163), .C2(new_n568), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1160), .A2(new_n1166), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1151), .A2(new_n1154), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1145), .A2(new_n1159), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1134), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1021), .A2(G286), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1107), .A2(new_n1118), .A3(new_n1119), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT116), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1098), .A2(new_n1180), .A3(new_n1107), .A4(new_n1177), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1107), .A2(KEYINPUT63), .A3(new_n1119), .A4(new_n1177), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1099), .B1(new_n1186), .B2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1184), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(G8), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1089), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1177), .A2(new_n1119), .A3(KEYINPUT63), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1190), .A2(KEYINPUT118), .A3(new_n1107), .A4(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1183), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1107), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1080), .A2(new_n1082), .A3(new_n834), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1078), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1194), .A2(new_n1119), .B1(new_n1076), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1122), .A2(new_n1176), .A3(new_n1193), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1050), .A2(new_n1017), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(G1996), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT111), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1199), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n884), .A2(G2067), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n789), .A2(new_n1156), .ZN(new_n1204));
  INV_X1    g779(.A(G1996), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n746), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1201), .A2(new_n746), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT112), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n896), .A2(new_n852), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n849), .A2(new_n851), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1202), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g789(.A(G290), .B(G1986), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1202), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1198), .A2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1201), .B(KEYINPUT46), .Z(new_n1218));
  INV_X1    g793(.A(KEYINPUT47), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1203), .A2(new_n746), .A3(new_n1204), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n1202), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1219), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n1199), .A2(G1986), .A3(G290), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1225), .B(KEYINPUT48), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1223), .A2(new_n1224), .B1(new_n1214), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1199), .B1(new_n1228), .B2(new_n1204), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1217), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1217), .A2(KEYINPUT126), .A3(new_n1230), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g810(.A1(G227), .A2(new_n459), .ZN(new_n1237));
  INV_X1    g811(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n675), .B2(new_n677), .ZN(new_n1239));
  OAI211_X1 g813(.A(new_n717), .B(new_n1239), .C1(new_n918), .C2(new_n920), .ZN(new_n1240));
  NOR3_X1   g814(.A1(new_n978), .A2(new_n976), .A3(new_n926), .ZN(new_n1241));
  OAI21_X1  g815(.A(KEYINPUT43), .B1(new_n1241), .B2(new_n974), .ZN(new_n1242));
  AOI211_X1 g816(.A(KEYINPUT127), .B(new_n1240), .C1(new_n1242), .C2(new_n999), .ZN(new_n1243));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1244));
  INV_X1    g818(.A(new_n1240), .ZN(new_n1245));
  AOI21_X1  g819(.A(new_n1244), .B1(new_n1000), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g820(.A1(new_n1243), .A2(new_n1246), .ZN(G308));
  NAND2_X1  g821(.A1(new_n1000), .A2(new_n1245), .ZN(G225));
endmodule


