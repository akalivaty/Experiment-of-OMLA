//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XNOR2_X1  g028(.A(G325), .B(KEYINPUT64), .ZN(G261));
  AND2_X1   g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n455), .A2(KEYINPUT65), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(KEYINPUT65), .B1(G567), .B2(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n467), .A2(new_n468), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n485), .B2(G138), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT67), .A2(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT67), .A2(G114), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n497), .B(G2105), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT67), .A2(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n465), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n497), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n500), .B(G2104), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  OAI21_X1  g084(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n475), .B1(new_n510), .B2(new_n506), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(new_n500), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n496), .B1(new_n509), .B2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n522), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  XNOR2_X1  g107(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n525), .A2(G51), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G89), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n535), .A2(new_n536), .A3(new_n539), .A4(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  AOI22_X1  g117(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n521), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n525), .A2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n517), .A2(new_n518), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n525), .A2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n528), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n552), .A2(KEYINPUT73), .A3(G651), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n537), .A2(G91), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n527), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n525), .A2(new_n574), .A3(G53), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n550), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n573), .A2(new_n575), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n570), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  AOI22_X1  g157(.A1(new_n537), .A2(G87), .B1(new_n525), .B2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  NAND3_X1  g160(.A1(new_n527), .A2(G48), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n525), .A2(KEYINPUT77), .A3(G48), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(new_n589), .B1(G86), .B2(new_n537), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n517), .B2(new_n518), .ZN(new_n592));
  AND2_X1   g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n537), .A2(G85), .B1(new_n525), .B2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n521), .B2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(KEYINPUT78), .B(G66), .Z(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n550), .A2(new_n604), .B1(new_n605), .B2(new_n516), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI221_X1 g183(.A(KEYINPUT79), .B1(new_n605), .B2(new_n516), .C1(new_n550), .C2(new_n604), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n608), .A2(G651), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n528), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(G54), .B2(new_n525), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n603), .B1(new_n618), .B2(new_n602), .ZN(G321));
  XOR2_X1   g194(.A(G321), .B(KEYINPUT81), .Z(G284));
  NAND2_X1  g195(.A1(G299), .A2(new_n602), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n618), .B1(new_n624), .B2(G860), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT82), .ZN(G148));
  NOR2_X1   g201(.A1(new_n563), .A2(G868), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n610), .A2(new_n615), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n616), .A2(KEYINPUT80), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n631), .B2(G868), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n463), .A2(new_n476), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT85), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n481), .A2(G123), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n485), .A2(G135), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n465), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n640), .A2(new_n642), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n638), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n648), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n684), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n688), .C1(new_n682), .C2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G2084), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(KEYINPUT24), .B2(G34), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n701));
  INV_X1    g276(.A(G160), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G33), .ZN(new_n704));
  NAND2_X1  g279(.A1(G115), .A2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(G127), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n480), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n465), .B1(new_n707), .B2(KEYINPUT94), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT94), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n710));
  NAND2_X1  g285(.A1(G103), .A2(G2104), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n485), .A2(G139), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n704), .B1(new_n715), .B2(new_n699), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n698), .A2(new_n703), .B1(new_n716), .B2(G2072), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n699), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n699), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT29), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n717), .B1(G2072), .B2(new_n716), .C1(new_n721), .C2(G2090), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n723), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n725), .A2(G1966), .B1(new_n727), .B2(G1961), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(G1961), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(G1966), .C2(new_n725), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT31), .B(G11), .Z(new_n731));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n699), .B1(new_n732), .B2(G28), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(KEYINPUT97), .B1(new_n732), .B2(G28), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n647), .B2(new_n699), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n699), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n481), .A2(G128), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n485), .A2(G140), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n699), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n739), .B1(G2067), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT98), .B2(new_n738), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n752), .C1(new_n703), .C2(new_n698), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n722), .A2(new_n730), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G164), .A2(new_n699), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G27), .B2(new_n699), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT99), .B(G2078), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n563), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G16), .B2(G19), .ZN(new_n760));
  INV_X1    g335(.A(G1341), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(new_n756), .B2(new_n757), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n758), .B(new_n762), .C1(new_n761), .C2(new_n760), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n699), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n481), .A2(G129), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n476), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n699), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n723), .A2(G20), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G2090), .B2(new_n721), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n776), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n777), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n723), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n618), .B2(new_n723), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT93), .B(G1348), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n764), .A2(new_n785), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n792));
  NOR2_X1   g367(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G6), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G305), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT90), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n723), .A2(G22), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G303), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n723), .A2(G23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G288), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n802), .A2(new_n804), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n802), .A2(new_n813), .A3(KEYINPUT34), .A4(new_n804), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  INV_X1    g395(.A(G1986), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n481), .A2(G119), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n485), .A2(G131), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n465), .A2(G107), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G25), .B(new_n828), .S(G29), .Z(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n822), .A2(new_n823), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n792), .B(new_n794), .C1(new_n818), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n816), .B2(new_n817), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT92), .B1(new_n834), .B2(new_n793), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n833), .A2(new_n841), .A3(new_n835), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n791), .B1(new_n840), .B2(new_n842), .ZN(G311));
  INV_X1    g418(.A(new_n791), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n841), .B1(new_n833), .B2(new_n835), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(G150));
  XNOR2_X1  g422(.A(KEYINPUT104), .B(G860), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n618), .A2(G559), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n521), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n525), .A2(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n528), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n560), .B2(new_n562), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n558), .B1(new_n553), .B2(new_n554), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n855), .A2(new_n858), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n561), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n853), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n849), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n862), .A2(new_n848), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n772), .B(new_n747), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n875), .B2(G2105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n485), .A2(G142), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT105), .Z(new_n878));
  AOI211_X1 g453(.A(new_n876), .B(new_n878), .C1(G130), .C2(new_n481), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n873), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n485), .A2(new_n492), .A3(G138), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n881), .A2(new_n882), .B1(new_n481), .B2(G126), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n512), .B1(new_n511), .B2(new_n500), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n715), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n828), .B(new_n636), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n880), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G160), .B(new_n647), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n890), .A2(new_n892), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(G395));
  XOR2_X1   g476(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n864), .A2(KEYINPUT107), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n860), .A2(new_n904), .A3(new_n863), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n903), .A2(new_n624), .A3(new_n618), .A4(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n860), .A2(new_n904), .A3(new_n863), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n860), .B2(new_n863), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n631), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n616), .A2(G299), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n616), .A2(G299), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n628), .A2(new_n570), .A3(new_n580), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n616), .A2(G299), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(KEYINPUT108), .A3(new_n914), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n906), .A2(new_n909), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n906), .A2(new_n909), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n902), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n906), .A2(new_n909), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n902), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n906), .A2(new_n909), .A3(new_n922), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G305), .B(G290), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n924), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n862), .A2(G868), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(G295));
  NOR3_X1   g516(.A1(new_n921), .A2(new_n923), .A3(new_n902), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n602), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n945), .B2(new_n939), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n938), .A2(new_n947), .A3(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(G171), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT112), .B1(new_n544), .B2(new_n547), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(G168), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(G301), .A2(KEYINPUT112), .A3(G286), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n865), .A2(new_n956), .A3(KEYINPUT114), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n860), .A2(new_n953), .A3(new_n863), .A4(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n864), .A2(new_n955), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n957), .A2(new_n919), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n865), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(KEYINPUT113), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n962), .B(new_n933), .C1(new_n967), .C2(new_n926), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n968), .A2(new_n894), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n962), .B1(new_n967), .B2(new_n926), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n934), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n912), .A2(new_n916), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n957), .A2(new_n961), .A3(new_n960), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n965), .A2(new_n966), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n963), .A2(new_n922), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n974), .A2(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n968), .B(new_n894), .C1(new_n978), .C2(new_n933), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n979), .B2(KEYINPUT43), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n973), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n970), .B1(new_n969), .B2(new_n972), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(G397));
  XNOR2_X1  g563(.A(new_n746), .B(new_n751), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT117), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n772), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n886), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n474), .A2(G40), .A3(new_n477), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n469), .A2(new_n461), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT66), .B1(new_n998), .B2(G2105), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n460), .B(new_n465), .C1(new_n469), .C2(new_n461), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT116), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n472), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n991), .A2(new_n993), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n992), .A3(new_n772), .ZN(new_n1008));
  INV_X1    g583(.A(new_n830), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n828), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n828), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  INV_X1    g591(.A(G1966), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n886), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1005), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1021), .B2(new_n995), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1002), .A2(new_n1004), .B1(new_n886), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT119), .B(G2084), .Z(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1016), .B(G8), .C1(new_n1028), .C2(G286), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1002), .A2(new_n1004), .B1(new_n886), .B2(new_n1019), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1018), .B1(G164), .B2(G1384), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1966), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G286), .A2(G8), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(KEYINPUT51), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT124), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1039), .B(new_n1035), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1029), .B(new_n1036), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n509), .A2(new_n513), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n1043), .B2(new_n883), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1003), .B1(new_n472), .B2(new_n997), .ZN(new_n1045));
  AOI211_X1 g620(.A(KEYINPUT116), .B(new_n996), .C1(new_n466), .C2(new_n471), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G288), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G1976), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1047), .A2(G8), .A3(new_n1049), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n590), .B(new_n1055), .C1(new_n596), .C2(new_n597), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n588), .A2(new_n589), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n537), .A2(G86), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n594), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(new_n1060), .A3(KEYINPUT49), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n1047), .A3(new_n1064), .A4(G8), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1051), .A2(new_n1054), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n1044), .B2(KEYINPUT45), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1069), .B(new_n1018), .C1(G164), .C2(G1384), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1031), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n807), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1024), .A2(new_n1073), .A3(new_n1025), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G303), .A2(G8), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT55), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1067), .B(new_n1077), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1068), .A2(new_n1031), .A3(new_n1070), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1023), .ZN(new_n1086));
  OAI22_X1  g661(.A1(new_n1045), .A2(new_n1046), .B1(G164), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT50), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1044), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1031), .A2(new_n1032), .A3(KEYINPUT53), .A4(new_n1081), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(G171), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1079), .A2(new_n1080), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1037), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1039), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1028), .A2(KEYINPUT124), .A3(new_n1037), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1036), .A4(new_n1029), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1042), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1047), .A2(G8), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1065), .A2(new_n1052), .A3(new_n1048), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1056), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1080), .B2(new_n1066), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT56), .B(G2072), .Z(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT121), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1068), .A2(new_n1031), .A3(new_n1070), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n782), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT120), .B1(new_n573), .B2(new_n575), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT57), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G299), .B(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1348), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1005), .A2(new_n751), .A3(new_n1044), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n628), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1068), .A2(new_n1031), .A3(new_n1070), .A4(new_n992), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1047), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT123), .B1(new_n1127), .B2(KEYINPUT59), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n563), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n563), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1128), .ZN(new_n1132));
  INV_X1    g707(.A(G1348), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1119), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n628), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1112), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1114), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT61), .B1(new_n1117), .B2(new_n1113), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1122), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NOR4_X1   g724(.A1(new_n996), .A2(new_n470), .A3(new_n1083), .A4(G2078), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1020), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(new_n995), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1032), .A2(KEYINPUT125), .A3(new_n1020), .A4(new_n1150), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1090), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1084), .A2(new_n1154), .A3(G171), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1157));
  AOI21_X1  g732(.A(G301), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1148), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(G171), .B1(new_n1084), .B2(new_n1154), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(G301), .A3(new_n1157), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(KEYINPUT54), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1147), .A2(new_n1159), .A3(new_n1041), .A4(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1101), .B(new_n1105), .C1(new_n1146), .C2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1080), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1034), .A2(G286), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1066), .A4(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT63), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1015), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1006), .A2(new_n992), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT46), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n991), .A2(new_n1006), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1011), .B(KEYINPUT126), .Z(new_n1176));
  NAND3_X1  g751(.A1(new_n1007), .A2(new_n1008), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(G2067), .B2(new_n746), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1006), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1006), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  OAI211_X1 g757(.A(new_n1175), .B(new_n1179), .C1(new_n1013), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g760(.A1(new_n458), .A2(G227), .ZN(new_n1187));
  AOI211_X1 g761(.A(G229), .B(new_n1187), .C1(new_n664), .C2(new_n666), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n895), .B2(new_n896), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1189), .A2(new_n986), .ZN(G308));
  OAI221_X1 g764(.A(new_n1188), .B1(new_n895), .B2(new_n896), .C1(new_n984), .C2(new_n985), .ZN(G225));
endmodule


