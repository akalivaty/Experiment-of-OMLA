

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608;

  XNOR2_X1 U327 ( .A(n397), .B(n396), .ZN(n558) );
  AND2_X1 U328 ( .A1(n393), .A2(n392), .ZN(n397) );
  BUF_X2 U329 ( .A(n561), .Z(n295) );
  XOR2_X1 U330 ( .A(n477), .B(n476), .Z(n561) );
  NOR2_X1 U331 ( .A1(n383), .A2(n388), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U333 ( .A(KEYINPUT99), .ZN(n409) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n462) );
  XOR2_X1 U335 ( .A(n424), .B(n364), .Z(n296) );
  XOR2_X1 U336 ( .A(KEYINPUT40), .B(n538), .Z(n297) );
  XOR2_X1 U337 ( .A(n465), .B(G99GAT), .Z(n298) );
  XOR2_X1 U338 ( .A(KEYINPUT30), .B(G8GAT), .Z(n299) );
  XNOR2_X1 U339 ( .A(n493), .B(KEYINPUT103), .ZN(n494) );
  NOR2_X1 U340 ( .A1(n558), .A2(n545), .ZN(n417) );
  XOR2_X1 U341 ( .A(G22GAT), .B(G155GAT), .Z(n447) );
  XOR2_X1 U342 ( .A(G8GAT), .B(G183GAT), .Z(n404) );
  XNOR2_X1 U343 ( .A(n308), .B(n307), .ZN(n313) );
  XNOR2_X1 U344 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U345 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U346 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U347 ( .A(n355), .B(KEYINPUT15), .ZN(n356) );
  NOR2_X1 U348 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U349 ( .A(n412), .B(n411), .ZN(n415) );
  XNOR2_X1 U350 ( .A(n357), .B(n356), .ZN(n358) );
  NOR2_X1 U351 ( .A1(n532), .A2(n541), .ZN(n509) );
  XOR2_X1 U352 ( .A(n471), .B(n470), .Z(n477) );
  XOR2_X1 U353 ( .A(n384), .B(KEYINPUT41), .Z(n578) );
  XOR2_X1 U354 ( .A(n381), .B(n380), .Z(n573) );
  INV_X1 U355 ( .A(G106GAT), .ZN(n513) );
  XNOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n483) );
  XNOR2_X1 U357 ( .A(n513), .B(KEYINPUT44), .ZN(n514) );
  XNOR2_X1 U358 ( .A(n510), .B(G92GAT), .ZN(n511) );
  XNOR2_X1 U359 ( .A(n515), .B(n514), .ZN(G1339GAT) );
  XNOR2_X1 U360 ( .A(n512), .B(n511), .ZN(G1337GAT) );
  XOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .Z(n301) );
  XNOR2_X1 U362 ( .A(G92GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n321) );
  INV_X1 U364 ( .A(G204GAT), .ZN(n302) );
  XNOR2_X1 U365 ( .A(n321), .B(n302), .ZN(n308) );
  XOR2_X1 U366 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n304) );
  XNOR2_X1 U367 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n306) );
  NAND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n305) );
  XOR2_X1 U370 ( .A(G78GAT), .B(KEYINPUT76), .Z(n310) );
  XNOR2_X1 U371 ( .A(G148GAT), .B(KEYINPUT75), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n310), .B(n309), .ZN(n451) );
  XNOR2_X1 U373 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n311), .B(KEYINPUT74), .ZN(n354) );
  XOR2_X1 U375 ( .A(n451), .B(n354), .Z(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n315) );
  INV_X1 U377 ( .A(n315), .ZN(n314) );
  NAND2_X1 U378 ( .A1(n314), .A2(n462), .ZN(n318) );
  INV_X1 U379 ( .A(n462), .ZN(n316) );
  NAND2_X1 U380 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND2_X1 U381 ( .A1(n318), .A2(n317), .ZN(n319) );
  XOR2_X1 U382 ( .A(G176GAT), .B(G64GAT), .Z(n405) );
  XNOR2_X1 U383 ( .A(n319), .B(n405), .ZN(n384) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n320), .B(G218GAT), .ZN(n413) );
  XOR2_X1 U386 ( .A(n321), .B(n413), .Z(n342) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G162GAT), .Z(n448) );
  INV_X1 U388 ( .A(KEYINPUT11), .ZN(n322) );
  NAND2_X1 U389 ( .A1(KEYINPUT10), .A2(n322), .ZN(n325) );
  INV_X1 U390 ( .A(KEYINPUT10), .ZN(n323) );
  NAND2_X1 U391 ( .A1(n323), .A2(KEYINPUT11), .ZN(n324) );
  NAND2_X1 U392 ( .A1(n325), .A2(n324), .ZN(n327) );
  XNOR2_X1 U393 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n326) );
  XNOR2_X1 U394 ( .A(n327), .B(n326), .ZN(n329) );
  INV_X1 U395 ( .A(n329), .ZN(n328) );
  NAND2_X1 U396 ( .A1(n448), .A2(n328), .ZN(n332) );
  INV_X1 U397 ( .A(n448), .ZN(n330) );
  NAND2_X1 U398 ( .A1(n330), .A2(n329), .ZN(n331) );
  NAND2_X1 U399 ( .A1(n332), .A2(n331), .ZN(n334) );
  NAND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n334), .B(n333), .ZN(n336) );
  INV_X1 U402 ( .A(KEYINPUT78), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U404 ( .A(G29GAT), .B(G43GAT), .Z(n338) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n367) );
  XNOR2_X1 U407 ( .A(n367), .B(KEYINPUT79), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n383) );
  INV_X1 U410 ( .A(KEYINPUT80), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n383), .B(n343), .ZN(n518) );
  INV_X1 U412 ( .A(n518), .ZN(n482) );
  XOR2_X1 U413 ( .A(KEYINPUT36), .B(n482), .Z(n605) );
  XOR2_X1 U414 ( .A(KEYINPUT81), .B(G64GAT), .Z(n345) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(G1GAT), .ZN(n344) );
  XNOR2_X1 U416 ( .A(n345), .B(n344), .ZN(n359) );
  XOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n347) );
  XNOR2_X1 U418 ( .A(G127GAT), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U419 ( .A(n347), .B(n346), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n404), .B(n447), .ZN(n349) );
  XOR2_X1 U421 ( .A(G71GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U422 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U423 ( .A(n351), .B(n350), .ZN(n353) );
  AND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U425 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U426 ( .A(n354), .B(KEYINPUT12), .Z(n355) );
  XOR2_X1 U427 ( .A(n359), .B(n358), .Z(n601) );
  INV_X1 U428 ( .A(n601), .ZN(n582) );
  NOR2_X1 U429 ( .A1(n605), .A2(n582), .ZN(n360) );
  XOR2_X1 U430 ( .A(KEYINPUT45), .B(n360), .Z(n361) );
  NOR2_X1 U431 ( .A1(n384), .A2(n361), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n362), .B(KEYINPUT116), .ZN(n382) );
  XOR2_X1 U433 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(G50GAT), .ZN(n363) );
  XNOR2_X1 U435 ( .A(n299), .B(n363), .ZN(n364) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n296), .B(n365), .ZN(n366) );
  XNOR2_X1 U438 ( .A(n366), .B(G141GAT), .ZN(n369) );
  XOR2_X1 U439 ( .A(n367), .B(G197GAT), .Z(n368) );
  XNOR2_X1 U440 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT73), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT67), .B(KEYINPUT72), .ZN(n370) );
  XOR2_X1 U443 ( .A(n371), .B(n370), .Z(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n381) );
  XOR2_X1 U445 ( .A(KEYINPUT29), .B(G15GAT), .Z(n375) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(KEYINPUT66), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U448 ( .A(G22GAT), .B(KEYINPUT71), .Z(n377) );
  XNOR2_X1 U449 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n379), .B(n378), .ZN(n380) );
  NAND2_X1 U452 ( .A1(n382), .A2(n573), .ZN(n393) );
  INV_X1 U453 ( .A(n573), .ZN(n596) );
  NAND2_X1 U454 ( .A1(n596), .A2(n578), .ZN(n386) );
  XOR2_X1 U455 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n385) );
  XNOR2_X1 U456 ( .A(n386), .B(n385), .ZN(n387) );
  NAND2_X1 U457 ( .A1(n387), .A2(n582), .ZN(n388) );
  OR2_X1 U458 ( .A1(KEYINPUT47), .A2(n389), .ZN(n391) );
  NAND2_X1 U459 ( .A1(KEYINPUT47), .A2(n389), .ZN(n390) );
  NAND2_X1 U460 ( .A1(n391), .A2(n390), .ZN(n392) );
  INV_X1 U461 ( .A(KEYINPUT48), .ZN(n395) );
  INV_X1 U462 ( .A(KEYINPUT64), .ZN(n394) );
  XOR2_X1 U463 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n399) );
  XNOR2_X1 U464 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U466 ( .A(KEYINPUT17), .B(n400), .Z(n475) );
  XOR2_X1 U467 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n402) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(G204GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U470 ( .A(G211GAT), .B(n403), .Z(n446) );
  XOR2_X1 U471 ( .A(KEYINPUT100), .B(n404), .Z(n407) );
  XNOR2_X1 U472 ( .A(n405), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U474 ( .A(n446), .B(n408), .Z(n412) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n413), .B(KEYINPUT98), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X2 U478 ( .A(n475), .B(n416), .ZN(n545) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT54), .ZN(n441) );
  XOR2_X1 U480 ( .A(G127GAT), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT84), .B(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U483 ( .A(KEYINPUT85), .B(n420), .Z(n466) );
  XOR2_X1 U484 ( .A(G57GAT), .B(G148GAT), .Z(n422) );
  XNOR2_X1 U485 ( .A(G120GAT), .B(G162GAT), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n423), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U488 ( .A(G29GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n466), .B(n427), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n429) );
  XNOR2_X1 U492 ( .A(KEYINPUT1), .B(KEYINPUT96), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(KEYINPUT6), .B(n430), .Z(n432) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U497 ( .A(n433), .B(KEYINPUT97), .Z(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n435) );
  XNOR2_X1 U499 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U501 ( .A(KEYINPUT3), .B(n436), .Z(n452) );
  XNOR2_X1 U502 ( .A(n452), .B(G155GAT), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n553) );
  NAND2_X1 U505 ( .A1(n441), .A2(n553), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n442), .B(KEYINPUT65), .ZN(n594) );
  XOR2_X1 U507 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n444) );
  XNOR2_X1 U508 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n443) );
  XNOR2_X1 U509 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n460) );
  XOR2_X1 U511 ( .A(n447), .B(G218GAT), .Z(n450) );
  XNOR2_X1 U512 ( .A(G106GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n454) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U517 ( .A(n456), .B(n455), .Z(n458) );
  NAND2_X1 U518 ( .A1(G228GAT), .A2(G233GAT), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n497) );
  NAND2_X1 U521 ( .A1(n594), .A2(n497), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT55), .ZN(n478) );
  XOR2_X1 U523 ( .A(KEYINPUT86), .B(n462), .Z(n464) );
  NAND2_X1 U524 ( .A1(G227GAT), .A2(G233GAT), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U526 ( .A(G43GAT), .B(n466), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n298), .B(n467), .ZN(n471) );
  XOR2_X1 U528 ( .A(G176GAT), .B(G190GAT), .Z(n469) );
  XNOR2_X1 U529 ( .A(G15GAT), .B(G113GAT), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n473) );
  XNOR2_X1 U532 ( .A(G183GAT), .B(KEYINPUT89), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U535 ( .A(n295), .ZN(n496) );
  NAND2_X1 U536 ( .A1(n478), .A2(n496), .ZN(n479) );
  XNOR2_X2 U537 ( .A(KEYINPUT123), .B(n479), .ZN(n589) );
  NAND2_X1 U538 ( .A1(n589), .A2(n596), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  NAND2_X1 U541 ( .A1(n589), .A2(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  NAND2_X1 U543 ( .A1(n589), .A2(n578), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(G176GAT), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1349GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT27), .B(n545), .Z(n499) );
  INV_X1 U548 ( .A(n499), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n553), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT101), .B(n489), .ZN(n557) );
  INV_X1 U551 ( .A(n557), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n497), .B(KEYINPUT28), .ZN(n559) );
  AND2_X1 U553 ( .A1(n295), .A2(n559), .ZN(n490) );
  NAND2_X1 U554 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT102), .ZN(n505) );
  NOR2_X1 U556 ( .A1(n295), .A2(n545), .ZN(n493) );
  NAND2_X1 U557 ( .A1(n494), .A2(n497), .ZN(n495) );
  XOR2_X1 U558 ( .A(KEYINPUT25), .B(n495), .Z(n501) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT26), .ZN(n595) );
  NAND2_X1 U560 ( .A1(n595), .A2(n499), .ZN(n500) );
  NAND2_X1 U561 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U562 ( .A1(n502), .A2(n553), .ZN(n503) );
  NAND2_X1 U563 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U564 ( .A(n506), .B(KEYINPUT105), .ZN(n522) );
  NOR2_X1 U565 ( .A1(n605), .A2(n522), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n582), .ZN(n508) );
  XOR2_X1 U567 ( .A(KEYINPUT37), .B(n508), .Z(n532) );
  NAND2_X1 U568 ( .A1(n573), .A2(n578), .ZN(n541) );
  XOR2_X1 U569 ( .A(KEYINPUT112), .B(n509), .Z(n555) );
  NOR2_X1 U570 ( .A1(n555), .A2(n545), .ZN(n512) );
  XNOR2_X1 U571 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n510) );
  NOR2_X1 U572 ( .A1(n555), .A2(n559), .ZN(n515) );
  XOR2_X1 U573 ( .A(KEYINPUT108), .B(KEYINPUT34), .Z(n517) );
  XNOR2_X1 U574 ( .A(G1GAT), .B(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U575 ( .A(n517), .B(n516), .ZN(n525) );
  XOR2_X1 U576 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n520) );
  NAND2_X1 U577 ( .A1(n601), .A2(n518), .ZN(n519) );
  XNOR2_X1 U578 ( .A(n520), .B(n519), .ZN(n521) );
  NOR2_X1 U579 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(n523), .Z(n542) );
  OR2_X1 U581 ( .A1(n573), .A2(n384), .ZN(n531) );
  OR2_X1 U582 ( .A1(n542), .A2(n531), .ZN(n529) );
  NOR2_X1 U583 ( .A1(n553), .A2(n529), .ZN(n524) );
  XOR2_X1 U584 ( .A(n525), .B(n524), .Z(G1324GAT) );
  NOR2_X1 U585 ( .A1(n545), .A2(n529), .ZN(n526) );
  XOR2_X1 U586 ( .A(G8GAT), .B(n526), .Z(G1325GAT) );
  NOR2_X1 U587 ( .A1(n295), .A2(n529), .ZN(n528) );
  XNOR2_X1 U588 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n528), .B(n527), .ZN(G1326GAT) );
  NOR2_X1 U590 ( .A1(n559), .A2(n529), .ZN(n530) );
  XOR2_X1 U591 ( .A(G22GAT), .B(n530), .Z(G1327GAT) );
  NOR2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U593 ( .A(KEYINPUT38), .B(KEYINPUT109), .ZN(n533) );
  XNOR2_X1 U594 ( .A(n534), .B(n533), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n553), .A2(n539), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n535), .B(KEYINPUT39), .ZN(n536) );
  XNOR2_X1 U597 ( .A(G29GAT), .B(n536), .ZN(G1328GAT) );
  NOR2_X1 U598 ( .A1(n539), .A2(n545), .ZN(n537) );
  XOR2_X1 U599 ( .A(G36GAT), .B(n537), .Z(G1329GAT) );
  NOR2_X1 U600 ( .A1(n539), .A2(n295), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G43GAT), .B(n297), .ZN(G1330GAT) );
  NOR2_X1 U602 ( .A1(n539), .A2(n559), .ZN(n540) );
  XOR2_X1 U603 ( .A(G50GAT), .B(n540), .Z(G1331GAT) );
  OR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n553), .A2(n549), .ZN(n543) );
  XOR2_X1 U606 ( .A(n543), .B(KEYINPUT42), .Z(n544) );
  XNOR2_X1 U607 ( .A(G57GAT), .B(n544), .ZN(G1332GAT) );
  NOR2_X1 U608 ( .A1(n545), .A2(n549), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT110), .B(n546), .Z(n547) );
  XNOR2_X1 U610 ( .A(G64GAT), .B(n547), .ZN(G1333GAT) );
  NOR2_X1 U611 ( .A1(n295), .A2(n549), .ZN(n548) );
  XOR2_X1 U612 ( .A(G71GAT), .B(n548), .Z(G1334GAT) );
  NOR2_X1 U613 ( .A1(n559), .A2(n549), .ZN(n551) );
  XNOR2_X1 U614 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G78GAT), .B(n552), .Z(G1335GAT) );
  NOR2_X1 U617 ( .A1(n553), .A2(n555), .ZN(n554) );
  XOR2_X1 U618 ( .A(G85GAT), .B(n554), .Z(G1336GAT) );
  NOR2_X1 U619 ( .A1(n555), .A2(n295), .ZN(n556) );
  XOR2_X1 U620 ( .A(G99GAT), .B(n556), .Z(G1338GAT) );
  XOR2_X1 U621 ( .A(G113GAT), .B(KEYINPUT117), .Z(n563) );
  NOR2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n572) );
  NAND2_X1 U623 ( .A1(n572), .A2(n559), .ZN(n560) );
  NOR2_X1 U624 ( .A1(n295), .A2(n560), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n569), .A2(n596), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(G1340GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n565) );
  NAND2_X1 U628 ( .A1(n569), .A2(n578), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G120GAT), .B(n566), .ZN(G1341GAT) );
  NAND2_X1 U631 ( .A1(n569), .A2(n601), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT50), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G127GAT), .B(n568), .ZN(G1342GAT) );
  XOR2_X1 U634 ( .A(G134GAT), .B(KEYINPUT51), .Z(n571) );
  NAND2_X1 U635 ( .A1(n569), .A2(n482), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1343GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n595), .ZN(n585) );
  NOR2_X1 U638 ( .A1(n573), .A2(n585), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1344GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n577) );
  XNOR2_X1 U642 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  INV_X1 U644 ( .A(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n579), .A2(n585), .ZN(n580) );
  XOR2_X1 U646 ( .A(n581), .B(n580), .Z(G1345GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1346GAT) );
  INV_X1 U650 ( .A(n383), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT122), .B(n587), .Z(n588) );
  XNOR2_X1 U653 ( .A(G162GAT), .B(n588), .ZN(G1347GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n601), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n592) );
  XNOR2_X1 U657 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U659 ( .A(KEYINPUT125), .B(n593), .Z(n598) );
  NAND2_X1 U660 ( .A1(n594), .A2(n595), .ZN(n604) );
  INV_X1 U661 ( .A(n604), .ZN(n602) );
  NAND2_X1 U662 ( .A1(n602), .A2(n596), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n598), .B(n597), .ZN(G1352GAT) );
  XOR2_X1 U664 ( .A(G204GAT), .B(KEYINPUT61), .Z(n600) );
  NAND2_X1 U665 ( .A1(n602), .A2(n384), .ZN(n599) );
  XNOR2_X1 U666 ( .A(n600), .B(n599), .ZN(G1353GAT) );
  NAND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U668 ( .A(n603), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U669 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U670 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n606) );
  XNOR2_X1 U671 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U672 ( .A(G218GAT), .B(n608), .ZN(G1355GAT) );
endmodule

