//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT68), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n209), .A3(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT68), .B(G120gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n204), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n202), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G113gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G120gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n203), .B1(new_n206), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT23), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n233), .B(KEYINPUT25), .C1(new_n234), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT64), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n232), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT65), .B1(new_n247), .B2(KEYINPUT25), .ZN(new_n248));
  AND2_X1   g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n227), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(new_n229), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n237), .B(new_n238), .C1(new_n234), .C2(KEYINPUT64), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n242), .A2(KEYINPUT64), .A3(new_n243), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n228), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n241), .B1(new_n248), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n236), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT28), .ZN(new_n263));
  OR3_X1    g062(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n231), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n259), .A2(new_n261), .A3(new_n267), .A4(new_n236), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n263), .A2(new_n266), .A3(new_n242), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n262), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n268), .A4(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n225), .B1(new_n258), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n242), .A2(new_n243), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(new_n246), .A3(new_n237), .A4(new_n238), .ZN(new_n282));
  AOI211_X1 g081(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n282), .C2(new_n233), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n240), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n210), .A2(new_n211), .ZN(new_n286));
  INV_X1    g085(.A(new_n206), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n214), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n204), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n223), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n271), .A2(new_n273), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n278), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT32), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G15gat), .B(G43gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n275), .A2(new_n293), .ZN(new_n302));
  INV_X1    g101(.A(new_n278), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT34), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n302), .A2(new_n303), .B1(KEYINPUT70), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n300), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n294), .B(KEYINPUT32), .C1(new_n296), .C2(new_n307), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n301), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n301), .B2(new_n308), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n309), .A2(new_n310), .B1(KEYINPUT70), .B2(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n301), .A2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n305), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n301), .A2(new_n306), .A3(new_n308), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G50gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n323));
  OAI21_X1  g122(.A(G218gat), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n326), .B2(new_n327), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT77), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G155gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT77), .B(G155gat), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT78), .B(KEYINPUT2), .C1(new_n344), .C2(new_n336), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G141gat), .B(G148gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G155gat), .B(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  OR2_X1    g156(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT71), .B(KEYINPUT22), .Z(new_n361));
  OAI21_X1  g160(.A(new_n327), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n328), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n329), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n351), .A2(new_n333), .A3(new_n354), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n321), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n356), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n365), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n349), .B1(new_n343), .B2(new_n345), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n371), .A2(KEYINPUT3), .A3(new_n353), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(KEYINPUT84), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n320), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n320), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT3), .B1(new_n365), .B2(new_n321), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n371), .A2(new_n353), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT85), .B1(new_n379), .B2(new_n367), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n356), .A2(new_n373), .A3(new_n381), .A4(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G22gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n375), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n375), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n319), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n375), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n319), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n383), .A3(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n392), .A3(new_n394), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n317), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n285), .A2(new_n269), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n321), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n248), .A2(new_n257), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n274), .B1(new_n403), .B2(new_n240), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n370), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT75), .ZN(new_n412));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n285), .B2(new_n292), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT73), .B(new_n401), .C1(new_n404), .C2(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n405), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n423), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT74), .B1(new_n423), .B2(new_n370), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n410), .B(new_n417), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n370), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT74), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n409), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n426), .B1(new_n431), .B2(new_n414), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT30), .B1(new_n431), .B2(new_n414), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n399), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n410), .B(new_n414), .C1(new_n424), .C2(new_n425), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n416), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n410), .B1(new_n424), .B2(new_n425), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n415), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT87), .A4(new_n426), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G57gat), .ZN(new_n442));
  INV_X1    g241(.A(G85gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT3), .B1(new_n371), .B2(new_n353), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n215), .B2(new_n224), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n290), .A2(new_n223), .A3(KEYINPUT79), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n366), .A2(new_n445), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n378), .A2(new_n452), .A3(new_n225), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n378), .B2(new_n225), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT81), .A3(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n454), .A2(new_n455), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n460), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT80), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n453), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n460), .A4(new_n449), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n378), .A2(new_n225), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n448), .A2(new_n447), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n378), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n444), .B(new_n463), .C1(new_n470), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n444), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n466), .B2(new_n469), .ZN(new_n478));
  INV_X1    g277(.A(new_n462), .ZN(new_n479));
  AOI211_X1 g278(.A(new_n450), .B(new_n479), .C1(new_n456), .C2(new_n458), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n476), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT6), .B(new_n477), .C1(new_n478), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n398), .A2(new_n434), .A3(new_n439), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n476), .A2(new_n481), .A3(KEYINPUT82), .A4(new_n482), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n484), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n432), .A2(new_n433), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n387), .A2(new_n392), .A3(new_n394), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n394), .B1(new_n387), .B2(new_n392), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n496), .A4(new_n317), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n488), .A2(KEYINPUT92), .B1(KEYINPUT35), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n317), .A2(new_n396), .A3(new_n397), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n485), .A2(new_n486), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n434), .A4(new_n439), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n434), .A2(new_n439), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n505));
  OR3_X1    g304(.A1(new_n459), .A2(new_n460), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n473), .A2(new_n461), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT39), .B(new_n507), .C1(new_n459), .C2(new_n460), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n444), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT40), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n511), .A2(new_n481), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n431), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n424), .A2(new_n425), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n410), .A2(new_n515), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n415), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT38), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n414), .A2(KEYINPUT38), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n437), .A2(new_n515), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n423), .A2(new_n525), .A3(new_n370), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n423), .B2(new_n370), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n515), .B1(new_n408), .B2(new_n370), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n523), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n483), .A2(new_n484), .A3(new_n435), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT90), .B(KEYINPUT38), .C1(new_n516), .C2(new_n519), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n522), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n534), .A3(new_n496), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n317), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n494), .B2(new_n495), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n396), .A2(KEYINPUT86), .A3(new_n397), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n492), .A2(new_n493), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n498), .A2(new_n503), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT11), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(new_n226), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G197gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT93), .Z(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G1gat), .B2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G43gat), .B(G50gat), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(G29gat), .B2(G36gat), .ZN(new_n564));
  NOR3_X1   g363(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(new_n564), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G29gat), .A2(G36gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n565), .B2(KEYINPUT94), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n563), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n557), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(KEYINPUT17), .A3(new_n573), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n576), .A2(new_n577), .B1(new_n574), .B2(new_n557), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT18), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n574), .B(new_n556), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n579), .B(KEYINPUT13), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n580), .A2(KEYINPUT18), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n550), .A2(new_n581), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n581), .A3(new_n585), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n549), .B(KEYINPUT12), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n544), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT96), .B(G57gat), .Z(new_n594));
  MUX2_X1   g393(.A(G57gat), .B(new_n594), .S(G64gat), .Z(new_n595));
  XOR2_X1   g394(.A(G71gat), .B(G78gat), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n596), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n595), .B(new_n602), .C1(new_n597), .C2(new_n601), .ZN(new_n603));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n596), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT98), .ZN(new_n608));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT99), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n557), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n611), .B(new_n613), .Z(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n574), .A2(new_n575), .ZN(new_n624));
  NAND2_X1  g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  AOI22_X1  g427(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n443), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G99gat), .B(G106gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(new_n577), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n574), .A2(new_n632), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n640), .B(new_n643), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n626), .A2(new_n631), .A3(new_n629), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n606), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n632), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n606), .A2(new_n633), .A3(new_n649), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n632), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  INV_X1    g458(.A(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT104), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n647), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n647), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G176gat), .ZN(new_n665));
  INV_X1    g464(.A(G204gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n655), .A2(new_n657), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n646), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n671), .B2(new_n663), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n645), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n593), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n492), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(G1gat), .Z(G1324gat));
  INV_X1    g476(.A(new_n504), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n682), .B(new_n683), .C1(new_n555), .C2(new_n679), .ZN(G1325gat));
  XNOR2_X1  g483(.A(new_n317), .B(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n317), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n675), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n539), .A2(new_n540), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n623), .ZN(new_n695));
  INV_X1    g494(.A(new_n644), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n669), .A2(new_n672), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n593), .A2(new_n695), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G29gat), .A3(new_n492), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n544), .B2(new_n644), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n487), .A2(new_n496), .A3(new_n317), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT92), .B1(new_n703), .B2(new_n504), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n704), .A2(new_n503), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n436), .A2(new_n426), .A3(new_n438), .ZN(new_n707));
  INV_X1    g506(.A(new_n484), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n483), .B2(new_n489), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n491), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n685), .B1(new_n691), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n496), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n504), .B2(new_n513), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n534), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT44), .B(new_n696), .C1(new_n706), .C2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n702), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n623), .A2(new_n592), .A3(new_n673), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n492), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n719), .ZN(G1328gat));
  NOR3_X1   g519(.A1(new_n698), .A2(G36gat), .A3(new_n678), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n718), .B2(new_n678), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  NOR3_X1   g523(.A1(new_n698), .A2(G43gat), .A3(new_n688), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT106), .ZN(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n718), .B2(new_n685), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G43gat), .B1(new_n718), .B2(new_n686), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g530(.A1(new_n698), .A2(G50gat), .A3(new_n691), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G50gat), .B1(new_n718), .B2(new_n496), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n716), .A2(new_n541), .A3(new_n717), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n732), .B1(new_n737), .B2(G50gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g538(.A1(new_n544), .A2(new_n591), .A3(new_n645), .A4(new_n697), .ZN(new_n740));
  INV_X1    g539(.A(new_n492), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT107), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n594), .ZN(G1332gat));
  AND2_X1   g543(.A1(new_n740), .A2(new_n504), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  INV_X1    g548(.A(new_n686), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n599), .B1(new_n740), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n688), .A2(G71gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n740), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n541), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n623), .A2(new_n591), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n697), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n716), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n492), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n535), .A2(new_n543), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n704), .A2(new_n503), .A3(new_n705), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n644), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n673), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n741), .A2(new_n443), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n702), .A2(new_n504), .A3(new_n715), .A4(new_n759), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT108), .Z(new_n773));
  NOR2_X1   g572(.A1(new_n678), .A2(G92gat), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n766), .A2(KEYINPUT109), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n544), .A2(new_n644), .A3(new_n758), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n766), .A2(KEYINPUT109), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n764), .B2(new_n757), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n673), .B(new_n774), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT110), .Z(new_n780));
  OAI21_X1  g579(.A(KEYINPUT52), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  INV_X1    g581(.A(new_n774), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n772), .B(new_n782), .C1(new_n768), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n760), .A2(new_n786), .A3(new_n686), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n317), .A3(new_n673), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n786), .ZN(G1338gat));
  NOR3_X1   g588(.A1(new_n697), .A2(new_n496), .A3(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n767), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n702), .A2(new_n712), .A3(new_n715), .A4(new_n759), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n702), .A2(new_n541), .A3(new_n715), .A4(new_n759), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n790), .B1(new_n776), .B2(new_n778), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n796), .B1(new_n800), .B2(KEYINPUT53), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT111), .B(new_n792), .C1(new_n798), .C2(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n795), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT112), .B(new_n795), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n646), .C1(new_n659), .C2(new_n660), .ZN(new_n809));
  INV_X1    g608(.A(new_n667), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT54), .B1(new_n670), .B2(new_n646), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(KEYINPUT55), .C1(new_n662), .C2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n668), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n658), .A2(new_n661), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n647), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n811), .B1(new_n662), .B2(new_n812), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n813), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(new_n591), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n582), .A2(new_n584), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT114), .Z(new_n826));
  NOR2_X1   g625(.A1(new_n578), .A2(new_n579), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n548), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n673), .A2(new_n587), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n696), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n587), .A2(new_n828), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n644), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n818), .A2(new_n832), .A3(new_n821), .A4(new_n823), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n695), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n674), .A2(new_n592), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n492), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n398), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n678), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n218), .A3(new_n591), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n836), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(KEYINPUT115), .A3(new_n691), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT115), .B1(new_n841), .B2(new_n691), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n504), .A2(new_n492), .A3(new_n688), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n591), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(KEYINPUT116), .A3(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n846), .B2(G113gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n845), .ZN(new_n850));
  OAI21_X1  g649(.A(G120gat), .B1(new_n850), .B2(new_n697), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n839), .A2(new_n213), .A3(new_n673), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n850), .B2(new_n695), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n221), .A3(new_n623), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n678), .A2(new_n696), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(G134gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n696), .A3(new_n845), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n861), .A2(new_n862), .A3(G134gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n861), .B2(G134gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(G1343gat));
  NAND3_X1  g664(.A1(new_n837), .A2(new_n712), .A3(new_n686), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n866), .A2(G141gat), .A3(new_n592), .A4(new_n504), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n697), .A2(new_n831), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n821), .A2(new_n591), .ZN(new_n869));
  INV_X1    g668(.A(new_n817), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT118), .B1(new_n871), .B2(new_n696), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n821), .A2(new_n591), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n829), .B1(new_n873), .B2(new_n817), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n644), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n833), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n877), .A2(new_n695), .B1(new_n592), .B2(new_n674), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n878), .B2(new_n691), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n496), .B1(new_n835), .B2(new_n836), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n537), .A2(new_n504), .A3(new_n492), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n879), .A2(new_n591), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n867), .B1(G141gat), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT119), .B1(new_n884), .B2(G141gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  AOI221_X4 g687(.A(new_n867), .B1(KEYINPUT119), .B2(new_n888), .C1(G141gat), .C2(new_n884), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n866), .A2(new_n504), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n673), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n697), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n892), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n881), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n833), .B1(new_n871), .B2(new_n696), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n695), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT57), .B(new_n691), .C1(new_n900), .C2(new_n836), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n673), .A3(new_n883), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n893), .B1(new_n896), .B2(new_n904), .ZN(G1345gat));
  INV_X1    g704(.A(new_n344), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n894), .B2(new_n695), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n344), .A3(new_n623), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT120), .ZN(G1346gat));
  NOR3_X1   g709(.A1(new_n866), .A2(G162gat), .A3(new_n857), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT121), .ZN(new_n912));
  OAI21_X1  g711(.A(G162gat), .B1(new_n894), .B2(new_n644), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1347gat));
  NAND2_X1  g713(.A1(new_n504), .A2(new_n492), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n688), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n844), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n592), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n915), .A2(new_n499), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n841), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n226), .A3(new_n591), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT122), .Z(new_n922));
  NAND2_X1  g721(.A1(new_n918), .A2(new_n922), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n917), .B2(new_n697), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n227), .A3(new_n673), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  AND2_X1   g725(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g726(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n259), .A2(new_n261), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n841), .A2(new_n929), .A3(new_n623), .A4(new_n919), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT123), .Z(new_n931));
  OAI211_X1 g730(.A(new_n623), .B(new_n916), .C1(new_n842), .C2(new_n843), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G183gat), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n927), .B(new_n928), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  AND4_X1   g733(.A1(KEYINPUT124), .A2(new_n931), .A3(new_n933), .A4(KEYINPUT60), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n236), .A3(new_n696), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n844), .A2(new_n696), .A3(new_n916), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(G190gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n938), .B2(G190gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n750), .A2(new_n915), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n880), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g743(.A(KEYINPUT125), .B(G197gat), .Z(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n591), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n902), .A2(new_n943), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n592), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n945), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n666), .A3(new_n673), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  AND3_X1   g750(.A1(new_n902), .A2(new_n673), .A3(new_n943), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n666), .B2(new_n952), .ZN(G1353gat));
  OAI21_X1  g752(.A(G211gat), .B1(new_n947), .B2(new_n695), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n944), .A2(new_n358), .A3(new_n359), .A4(new_n623), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n944), .B2(new_n696), .ZN(new_n960));
  INV_X1    g759(.A(new_n947), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n696), .A2(G218gat), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT127), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(G1355gat));
endmodule


