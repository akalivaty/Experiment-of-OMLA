//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT40), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT39), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G141gat), .B(G148gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT81), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n206), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G127gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G134gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT70), .B(G134gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(new_n222), .ZN(new_n225));
  XOR2_X1   g024(.A(G113gat), .B(G120gat), .Z(new_n226));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G134gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT1), .B1(new_n229), .B2(G127gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(G113gat), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n230), .A2(new_n233), .A3(new_n223), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT71), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n225), .A2(new_n228), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n221), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n220), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n214), .B2(new_n216), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n217), .A2(new_n247), .A3(new_n237), .A4(new_n220), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(KEYINPUT82), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n248), .B2(KEYINPUT82), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(new_n247), .B2(new_n239), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(KEYINPUT82), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT83), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n247), .B1(new_n241), .B2(new_n237), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(KEYINPUT82), .A3(new_n249), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n241), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n258), .A2(new_n237), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n252), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n203), .B(new_n246), .C1(new_n263), .C2(new_n245), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n203), .A3(new_n245), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  INV_X1    g065(.A(G85gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G57gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n264), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n245), .ZN(new_n274));
  INV_X1    g073(.A(new_n246), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT39), .A3(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(KEYINPUT40), .A3(new_n271), .A4(new_n265), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT65), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n289), .A2(G169gat), .A3(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n282), .A2(new_n285), .A3(new_n296), .A4(new_n286), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n281), .B1(new_n280), .B2(KEYINPUT66), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n280), .A2(KEYINPUT66), .A3(new_n281), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n284), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G190gat), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n302), .B(new_n303), .C1(new_n307), .C2(G183gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT25), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(G183gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n283), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(G183gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n311), .B1(new_n317), .B2(new_n307), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n311), .B1(new_n304), .B2(new_n306), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n291), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n291), .A2(new_n324), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT69), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n325), .A2(new_n293), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n322), .A2(new_n280), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n279), .B1(new_n310), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n306), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n301), .B1(new_n333), .B2(new_n283), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n334), .B2(new_n303), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n295), .A2(new_n335), .B1(new_n298), .B2(new_n299), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n315), .A3(new_n316), .A4(new_n314), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n337), .A2(new_n311), .B1(new_n320), .B2(new_n319), .ZN(new_n338));
  INV_X1    g137(.A(new_n280), .ZN(new_n339));
  INV_X1    g138(.A(new_n328), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n331), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n330), .B1(new_n342), .B2(new_n279), .ZN(new_n343));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(KEYINPUT22), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT74), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n343), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n348), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT74), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT29), .B1(new_n310), .B2(new_n329), .ZN(new_n357));
  INV_X1    g156(.A(new_n279), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n353), .B(new_n356), .C1(new_n359), .C2(new_n330), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n355), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT76), .B(G8gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(G36gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND4_X1  g164(.A1(new_n352), .A2(new_n360), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(KEYINPUT79), .A3(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n352), .A2(new_n361), .A3(new_n360), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT30), .A4(new_n365), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT78), .B1(new_n366), .B2(new_n367), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n352), .A2(new_n361), .A3(new_n360), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n365), .B(KEYINPUT77), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n252), .A2(new_n257), .A3(new_n262), .A4(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n245), .B1(new_n239), .B2(new_n242), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n255), .A2(new_n244), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n385), .A2(new_n248), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT5), .B(new_n384), .C1(new_n386), .C2(new_n261), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n271), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n278), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n358), .B1(new_n336), .B2(new_n341), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n391), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n392), .B(KEYINPUT37), .C1(new_n343), .C2(new_n350), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT88), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n355), .B1(new_n359), .B2(new_n330), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT37), .A4(new_n392), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n352), .A2(new_n360), .A3(new_n400), .A4(new_n361), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n379), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n378), .A2(KEYINPUT37), .ZN(new_n404));
  INV_X1    g203(.A(new_n365), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n401), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n402), .A2(new_n403), .B1(new_n406), .B2(KEYINPUT38), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n388), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT85), .B1(new_n388), .B2(KEYINPUT6), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT38), .B1(new_n394), .B2(new_n397), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n412), .A2(KEYINPUT89), .A3(new_n379), .A4(new_n401), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n383), .A2(new_n387), .A3(new_n271), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n416), .A2(new_n389), .B1(new_n373), .B2(new_n365), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n407), .A2(new_n411), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT31), .B(G50gat), .Z(new_n419));
  OAI21_X1  g218(.A(new_n331), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n350), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  INV_X1    g221(.A(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n259), .B1(new_n350), .B2(KEYINPUT29), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n221), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n356), .A2(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n419), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n429), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G22gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT86), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n440), .A3(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n390), .A2(new_n418), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(KEYINPUT87), .A3(new_n443), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n414), .A2(new_n450), .A3(new_n415), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n389), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n414), .B2(new_n415), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n410), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n408), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n449), .B1(new_n457), .B2(new_n381), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT72), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n238), .B1(new_n336), .B2(new_n341), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n310), .A2(new_n237), .A3(new_n329), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT72), .B(new_n463), .C1(new_n460), .C2(new_n461), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT32), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n463), .A3(new_n461), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n463), .B2(KEYINPUT73), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n460), .A2(new_n463), .A3(new_n461), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G43gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n310), .A2(new_n237), .A3(new_n329), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n237), .B1(new_n310), .B2(new_n329), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n464), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT72), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n459), .A3(new_n464), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n473), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(KEYINPUT32), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n475), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n486), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n475), .A2(new_n489), .B1(new_n491), .B2(new_n478), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT36), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n445), .A2(new_n458), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n490), .B2(new_n492), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n478), .ZN(new_n498));
  INV_X1    g297(.A(new_n489), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n488), .B1(new_n485), .B2(KEYINPUT32), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n475), .A2(new_n487), .A3(new_n489), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT90), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n375), .A2(new_n376), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n366), .A2(KEYINPUT79), .A3(new_n367), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT79), .B1(new_n366), .B2(new_n367), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n380), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n416), .A2(new_n389), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n455), .A3(new_n408), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n509), .A3(new_n444), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n452), .A2(new_n453), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n381), .B1(new_n514), .B2(new_n411), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n493), .A2(KEYINPUT35), .A3(new_n444), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n512), .A2(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G64gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G57gat), .ZN(new_n520));
  INV_X1    g319(.A(G57gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G64gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n525));
  INV_X1    g324(.A(G71gat), .ZN(new_n526));
  INV_X1    g325(.A(G78gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n525), .A3(new_n529), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n523), .A2(KEYINPUT9), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n528), .A2(new_n529), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n534), .B1(new_n520), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT96), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n533), .A2(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT21), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G8gat), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n544), .A2(new_n553), .A3(new_n283), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n283), .B1(new_n544), .B2(new_n553), .ZN(new_n555));
  INV_X1    g354(.A(G231gat), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n423), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n544), .A2(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G183gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n553), .A3(new_n283), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n556), .A2(new_n423), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n557), .B2(new_n562), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g367(.A(G211gat), .B1(new_n543), .B2(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n540), .A2(new_n542), .ZN(new_n570));
  INV_X1    g369(.A(new_n532), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n523), .B(new_n535), .C1(new_n571), .C2(new_n530), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT21), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n345), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n568), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n569), .A2(new_n575), .A3(new_n568), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n577), .B2(new_n580), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n566), .A2(new_n567), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n557), .A2(new_n562), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n563), .ZN(new_n586));
  INV_X1    g385(.A(new_n583), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n581), .A4(new_n565), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n267), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n267), .B2(new_n596), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT14), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT14), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(new_n609), .C1(G29gat), .C2(G36gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G29gat), .A2(G36gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(G29gat), .A2(G36gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n606), .A3(KEYINPUT14), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G43gat), .B(G50gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT15), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(KEYINPUT15), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n614), .B(new_n617), .C1(KEYINPUT92), .C2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n610), .A2(KEYINPUT92), .A3(new_n611), .A4(new_n613), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(new_n618), .C1(new_n622), .C2(new_n616), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(KEYINPUT100), .B2(new_n590), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n620), .B2(new_n623), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n620), .A2(new_n623), .A3(KEYINPUT93), .A4(new_n626), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n601), .B(new_n602), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n625), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n594), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND3_X1  g439(.A1(new_n634), .A2(new_n594), .A3(new_n635), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n636), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n589), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n518), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n631), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n550), .A2(new_n552), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT94), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n620), .A2(new_n623), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n648), .B(new_n650), .C1(new_n626), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n651), .B(new_n649), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n652), .A2(KEYINPUT18), .A3(new_n653), .A4(new_n654), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  INV_X1    g463(.A(G197gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT12), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n657), .A2(new_n661), .A3(new_n662), .A4(new_n669), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n543), .B2(new_n605), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT101), .B1(new_n543), .B2(new_n605), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n573), .A2(new_n677), .A3(new_n633), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n573), .B2(new_n633), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n543), .A2(new_n605), .A3(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n675), .B1(new_n684), .B2(new_n674), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n686), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT10), .B1(new_n679), .B2(new_n683), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n691), .A2(new_n692), .A3(new_n689), .A4(new_n675), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n688), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G120gat), .B(G148gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT104), .ZN(new_n697));
  XNOR2_X1  g496(.A(G176gat), .B(G204gat), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n697), .B(new_n698), .Z(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n686), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n699), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n673), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n647), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n457), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n381), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT16), .B(G8gat), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(G8gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n715), .A2(KEYINPUT106), .A3(new_n716), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1325gat));
  INV_X1    g521(.A(new_n494), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n709), .A2(G15gat), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(G15gat), .B1(new_n709), .B2(new_n504), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(G1326gat));
  INV_X1    g525(.A(new_n449), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NAND2_X1  g529(.A1(new_n645), .A2(new_n642), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n518), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n589), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n707), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n457), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(G29gat), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n645), .A2(new_n642), .A3(KEYINPUT108), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT108), .B1(new_n645), .B2(new_n642), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n518), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n518), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n741), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n734), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G29gat), .B1(new_n753), .B2(new_n737), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n754), .ZN(G1328gat));
  NOR3_X1   g554(.A1(new_n736), .A2(G36gat), .A3(new_n509), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g556(.A(G36gat), .B1(new_n753), .B2(new_n509), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1329gat));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  INV_X1    g559(.A(new_n731), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n495), .B2(new_n517), .ZN(new_n762));
  INV_X1    g561(.A(G43gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n763), .A3(new_n752), .ZN(new_n764));
  INV_X1    g563(.A(new_n504), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n764), .A2(KEYINPUT111), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT111), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n723), .A3(new_n752), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(G43gat), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(G43gat), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT110), .B(KEYINPUT47), .C1(new_n773), .C2(new_n768), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(G1330gat));
  AOI21_X1  g574(.A(new_n727), .B1(new_n736), .B2(KEYINPUT112), .ZN(new_n776));
  INV_X1    g575(.A(G50gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n776), .B(new_n777), .C1(KEYINPUT112), .C2(new_n736), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n753), .A2(new_n727), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n777), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G50gat), .B1(new_n753), .B2(new_n444), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n783), .A3(KEYINPUT48), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n778), .A2(new_n783), .A3(KEYINPUT113), .A4(KEYINPUT48), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(G1331gat));
  NAND4_X1  g587(.A1(new_n518), .A2(new_n673), .A3(new_n706), .A4(new_n646), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n737), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(new_n521), .ZN(G1332gat));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n381), .A3(new_n791), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT49), .B(G64gat), .Z(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(G1333gat));
  OAI21_X1  g597(.A(new_n526), .B1(new_n792), .B2(new_n765), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n790), .A2(G71gat), .A3(new_n723), .A4(new_n791), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n799), .B(new_n804), .C1(new_n801), .C2(new_n802), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1334gat));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n727), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(new_n527), .ZN(G1335gat));
  INV_X1    g609(.A(new_n705), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n695), .B2(new_n700), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n671), .A2(new_n672), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n589), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n751), .A2(KEYINPUT117), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT117), .B1(new_n751), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n457), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n457), .C1(new_n815), .C2(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(G85gat), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n813), .A2(new_n589), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n762), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n762), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n706), .A3(new_n826), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n827), .A2(G85gat), .A3(new_n737), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n828), .ZN(G1336gat));
  NOR3_X1   g628(.A1(new_n827), .A2(G92gat), .A3(new_n509), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n751), .A2(new_n814), .ZN(new_n832));
  OAI21_X1  g631(.A(G92gat), .B1(new_n832), .B2(new_n509), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n381), .B1(new_n815), .B2(new_n816), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n830), .B1(new_n835), .B2(G92gat), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(G1337gat));
  NOR2_X1   g637(.A1(new_n815), .A2(new_n816), .ZN(new_n839));
  OAI21_X1  g638(.A(G99gat), .B1(new_n839), .B2(new_n494), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n827), .A2(G99gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n765), .B2(new_n841), .ZN(G1338gat));
  OAI21_X1  g641(.A(G106gat), .B1(new_n832), .B2(new_n444), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n444), .A2(G106gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n843), .A2(new_n846), .A3(new_n850), .A4(new_n847), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n449), .B1(new_n815), .B2(new_n816), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n845), .B1(new_n852), .B2(G106gat), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n849), .B(new_n851), .C1(new_n853), .C2(new_n847), .ZN(G1339gat));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n731), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n742), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n687), .B2(new_n693), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n689), .B1(new_n691), .B2(new_n675), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n703), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n700), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n700), .A4(new_n861), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(new_n813), .A3(new_n705), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n654), .B1(new_n652), .B2(new_n653), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n658), .A2(new_n660), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n668), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n672), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n706), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n857), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n864), .A2(new_n705), .A3(new_n870), .A4(new_n865), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n745), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n733), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n646), .A2(new_n673), .A3(new_n812), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n646), .A2(new_n673), .A3(KEYINPUT120), .A4(new_n812), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n727), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n765), .B1(new_n882), .B2(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n457), .A2(new_n509), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n886), .A3(new_n727), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G113gat), .B1(new_n888), .B2(new_n673), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n881), .A2(new_n493), .A3(new_n444), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n885), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n891), .A2(G113gat), .A3(new_n673), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n888), .B2(new_n812), .ZN(new_n894));
  INV_X1    g693(.A(new_n891), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n232), .A3(new_n706), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1341gat));
  NOR3_X1   g696(.A1(new_n888), .A2(new_n222), .A3(new_n733), .ZN(new_n898));
  AOI21_X1  g697(.A(G127gat), .B1(new_n895), .B2(new_n589), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1342gat));
  NOR3_X1   g699(.A1(new_n891), .A2(new_n224), .A3(new_n761), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT56), .ZN(new_n902));
  OAI21_X1  g701(.A(G134gat), .B1(new_n888), .B2(new_n761), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1343gat));
  XNOR2_X1  g703(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n878), .A2(new_n879), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n866), .A2(new_n871), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n745), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n745), .A2(new_n873), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(new_n733), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT123), .B(new_n906), .C1(new_n912), .C2(new_n444), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n444), .B1(new_n875), .B2(new_n880), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n905), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n731), .B1(new_n866), .B2(new_n871), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n874), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n880), .B1(new_n918), .B2(new_n589), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(KEYINPUT57), .A3(new_n449), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n913), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n723), .A2(new_n884), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G141gat), .B1(new_n923), .B2(new_n673), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n915), .A2(new_n922), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n813), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(G141gat), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g727(.A(KEYINPUT124), .B(KEYINPUT58), .Z(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1344gat));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n706), .A3(new_n922), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(G148gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n912), .A2(new_n444), .A3(new_n906), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n873), .A2(new_n761), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n733), .B1(new_n917), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n876), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT57), .B1(new_n937), .B2(new_n449), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n922), .B(new_n706), .C1(new_n934), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G148gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n925), .A2(G148gat), .A3(new_n812), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1345gat));
  AOI21_X1  g747(.A(G155gat), .B1(new_n926), .B2(new_n589), .ZN(new_n949));
  INV_X1    g748(.A(new_n923), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n589), .A2(G155gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(G1346gat));
  AOI21_X1  g751(.A(G162gat), .B1(new_n926), .B2(new_n731), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n923), .A2(new_n745), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n457), .A2(new_n509), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n890), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(G169gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n813), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n961), .A2(new_n504), .A3(new_n887), .A4(new_n956), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n883), .A2(KEYINPUT126), .A3(new_n887), .A4(new_n956), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n964), .A2(new_n813), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n960), .B1(new_n966), .B2(new_n959), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n958), .B2(new_n706), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n964), .A2(new_n706), .A3(new_n965), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n589), .A3(new_n965), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G183gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n320), .A3(new_n589), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT60), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n958), .A2(new_n333), .A3(new_n857), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n731), .A3(new_n965), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n980), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n980), .B2(G190gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1351gat));
  NOR3_X1   g783(.A1(new_n723), .A2(new_n509), .A3(new_n444), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n912), .A2(new_n457), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n665), .A3(new_n813), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n934), .A2(new_n938), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(new_n494), .A3(new_n956), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(new_n813), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n994), .B2(new_n665), .ZN(G1352gat));
  NOR3_X1   g794(.A1(new_n988), .A2(G204gat), .A3(new_n812), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n996), .B(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n991), .A2(new_n706), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n956), .A2(new_n494), .ZN(new_n999));
  OAI21_X1  g798(.A(G204gat), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n997), .A2(new_n1000), .ZN(G1353gat));
  NAND3_X1  g800(.A1(new_n989), .A2(new_n345), .A3(new_n589), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n992), .A2(new_n589), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n346), .A3(new_n857), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n731), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1007), .B1(new_n1009), .B2(new_n346), .ZN(G1355gat));
endmodule


