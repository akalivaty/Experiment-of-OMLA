

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n755) );
  AND2_X2 U556 ( .A1(n530), .A2(G2104), .ZN(n878) );
  XOR2_X1 U557 ( .A(KEYINPUT93), .B(n689), .Z(n799) );
  XNOR2_X1 U558 ( .A(n740), .B(n739), .ZN(n796) );
  OR2_X1 U559 ( .A1(n796), .A2(n795), .ZN(n806) );
  NAND2_X1 U560 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U561 ( .A(n524), .B(KEYINPUT65), .ZN(n519) );
  NOR2_X1 U562 ( .A1(n731), .A2(n947), .ZN(n698) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n702) );
  XNOR2_X1 U564 ( .A(n703), .B(n702), .ZN(n710) );
  XNOR2_X1 U565 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n695) );
  XNOR2_X1 U566 ( .A(n696), .B(n695), .ZN(n728) );
  INV_X1 U567 ( .A(n981), .ZN(n749) );
  NOR2_X1 U568 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X2 U569 ( .A1(G2104), .A2(n530), .ZN(n882) );
  NOR2_X1 U570 ( .A1(G651), .A2(n641), .ZN(n645) );
  NOR2_X1 U571 ( .A1(n641), .A2(n543), .ZN(n653) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n646) );
  NOR2_X2 U573 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U574 ( .A(G2105), .ZN(n530) );
  AND2_X1 U575 ( .A1(G2104), .A2(G101), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n530), .A2(n520), .ZN(n521) );
  XOR2_X1 U577 ( .A(n521), .B(KEYINPUT23), .Z(n523) );
  NAND2_X1 U578 ( .A1(n882), .A2(G125), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XOR2_X1 U581 ( .A(KEYINPUT17), .B(n525), .Z(n532) );
  BUF_X1 U582 ( .A(n532), .Z(n879) );
  NAND2_X1 U583 ( .A1(G137), .A2(n879), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n519), .A2(n526), .ZN(n529) );
  AND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U586 ( .A1(n883), .A2(G113), .ZN(n527) );
  XOR2_X1 U587 ( .A(KEYINPUT66), .B(n527), .Z(n528) );
  NAND2_X1 U588 ( .A1(n878), .A2(G102), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n531), .B(KEYINPUT88), .ZN(n534) );
  NAND2_X1 U590 ( .A1(G138), .A2(n532), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n535), .B(KEYINPUT89), .ZN(n540) );
  AND2_X1 U593 ( .A1(G114), .A2(n883), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G126), .A2(n882), .ZN(n536) );
  XNOR2_X1 U595 ( .A(KEYINPUT87), .B(n536), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(G164) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G69), .ZN(G235) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  NAND2_X1 U602 ( .A1(n646), .A2(G88), .ZN(n542) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(G651), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G75), .A2(n653), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G50), .A2(n645), .ZN(n547) );
  NOR2_X1 U608 ( .A1(G543), .A2(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT68), .B(KEYINPUT1), .Z(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n649) );
  NAND2_X1 U611 ( .A1(G62), .A2(n649), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(G166) );
  NAND2_X1 U614 ( .A1(G51), .A2(n645), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G63), .A2(n649), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n552), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n646), .A2(G89), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G76), .A2(n653), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(n556), .B(KEYINPUT5), .Z(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT74), .B(n559), .Z(n560) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  XNOR2_X1 U626 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G168), .ZN(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n828) );
  NAND2_X1 U631 ( .A1(n828), .A2(G567), .ZN(n563) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U633 ( .A1(G56), .A2(n649), .ZN(n564) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n564), .Z(n571) );
  NAND2_X1 U635 ( .A1(n646), .A2(G81), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT12), .B(n565), .Z(n568) );
  NAND2_X1 U637 ( .A1(G68), .A2(n653), .ZN(n566) );
  XOR2_X1 U638 ( .A(KEYINPUT72), .B(n566), .Z(n567) );
  XNOR2_X1 U639 ( .A(n569), .B(KEYINPUT13), .ZN(n570) );
  NOR2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n645), .A2(G43), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n989) );
  INV_X1 U643 ( .A(n989), .ZN(n574) );
  XOR2_X1 U644 ( .A(G860), .B(KEYINPUT73), .Z(n602) );
  NAND2_X1 U645 ( .A1(n574), .A2(n602), .ZN(G153) );
  NAND2_X1 U646 ( .A1(n646), .A2(G90), .ZN(n576) );
  NAND2_X1 U647 ( .A1(G77), .A2(n653), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U649 ( .A(KEYINPUT9), .B(n577), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n645), .A2(G52), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G64), .A2(n649), .ZN(n578) );
  AND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n649), .A2(G66), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G79), .A2(n653), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G54), .A2(n645), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G92), .A2(n646), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n588), .Z(n621) );
  INV_X1 U663 ( .A(n621), .ZN(n977) );
  INV_X1 U664 ( .A(G868), .ZN(n665) );
  NAND2_X1 U665 ( .A1(n977), .A2(n665), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U667 ( .A1(n649), .A2(G65), .ZN(n592) );
  NAND2_X1 U668 ( .A1(G78), .A2(n653), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n645), .A2(G53), .ZN(n593) );
  XOR2_X1 U671 ( .A(KEYINPUT70), .B(n593), .Z(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n646), .A2(G91), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT76), .ZN(n600) );
  NOR2_X1 U677 ( .A1(G286), .A2(n665), .ZN(n599) );
  NOR2_X1 U678 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U679 ( .A(G559), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n977), .A2(n603), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT16), .B(n604), .Z(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n989), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G868), .A2(n621), .ZN(n605) );
  NOR2_X1 U685 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U687 ( .A(KEYINPUT77), .B(n608), .Z(G282) );
  XOR2_X1 U688 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n610) );
  NAND2_X1 U689 ( .A1(G123), .A2(n882), .ZN(n609) );
  XNOR2_X1 U690 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT78), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n878), .A2(G99), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G135), .A2(n879), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G111), .A2(n883), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n919) );
  XNOR2_X1 U698 ( .A(n919), .B(G2096), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT80), .ZN(n620) );
  INV_X1 U700 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U702 ( .A1(n621), .A2(G559), .ZN(n662) );
  XNOR2_X1 U703 ( .A(n989), .B(n662), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n622), .A2(G860), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n649), .A2(G67), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G80), .A2(n653), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G55), .A2(n645), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G93), .A2(n646), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n664) );
  XOR2_X1 U712 ( .A(n629), .B(n664), .Z(G145) );
  XOR2_X1 U713 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n631) );
  NAND2_X1 U714 ( .A1(G73), .A2(n653), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n631), .B(n630), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G48), .A2(n645), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G86), .A2(n646), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n649), .A2(G61), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n645), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U725 ( .A1(n649), .A2(n640), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G87), .A2(n641), .ZN(n642) );
  XOR2_X1 U727 ( .A(KEYINPUT81), .B(n642), .Z(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G47), .A2(n645), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G85), .A2(n646), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G60), .A2(n649), .ZN(n650) );
  XNOR2_X1 U733 ( .A(KEYINPUT69), .B(n650), .ZN(n651) );
  NOR2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G72), .A2(n653), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(G290) );
  INV_X1 U737 ( .A(G299), .ZN(n971) );
  XNOR2_X1 U738 ( .A(G166), .B(n971), .ZN(n660) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(G305), .ZN(n656) );
  XNOR2_X1 U740 ( .A(n656), .B(G288), .ZN(n657) );
  XOR2_X1 U741 ( .A(n664), .B(n657), .Z(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(G290), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n989), .B(n661), .ZN(n897) );
  XNOR2_X1 U745 ( .A(n662), .B(n897), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G237), .A2(G235), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G120), .A2(n672), .ZN(n673) );
  XNOR2_X1 U758 ( .A(KEYINPUT85), .B(n673), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(G108), .ZN(n833) );
  NAND2_X1 U760 ( .A1(n833), .A2(G567), .ZN(n681) );
  NOR2_X1 U761 ( .A1(G219), .A2(G220), .ZN(n676) );
  XNOR2_X1 U762 ( .A(KEYINPUT22), .B(KEYINPUT83), .ZN(n675) );
  XNOR2_X1 U763 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n677), .A2(G218), .ZN(n678) );
  NAND2_X1 U765 ( .A1(G96), .A2(n678), .ZN(n832) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n832), .ZN(n679) );
  XNOR2_X1 U767 ( .A(KEYINPUT84), .B(n679), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n834) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n834), .A2(n682), .ZN(n831) );
  NAND2_X1 U771 ( .A1(n831), .A2(G36), .ZN(n683) );
  XNOR2_X1 U772 ( .A(KEYINPUT86), .B(n683), .ZN(G176) );
  INV_X1 U773 ( .A(G166), .ZN(G303) );
  XOR2_X1 U774 ( .A(G2078), .B(KEYINPUT25), .Z(n949) );
  INV_X1 U775 ( .A(n755), .ZN(n685) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n754) );
  NOR2_X1 U777 ( .A1(n685), .A2(n754), .ZN(n686) );
  INV_X1 U778 ( .A(n686), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n949), .A2(n731), .ZN(n688) );
  BUF_X1 U780 ( .A(n686), .Z(n714) );
  XNOR2_X1 U781 ( .A(G1961), .B(KEYINPUT94), .ZN(n1014) );
  NOR2_X1 U782 ( .A1(n714), .A2(n1014), .ZN(n687) );
  NOR2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n724) );
  AND2_X1 U784 ( .A1(G301), .A2(n724), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n731), .A2(G8), .ZN(n689) );
  NOR2_X1 U786 ( .A1(G1966), .A2(n799), .ZN(n744) );
  NOR2_X1 U787 ( .A1(G2084), .A2(n731), .ZN(n741) );
  NOR2_X1 U788 ( .A1(n744), .A2(n741), .ZN(n690) );
  NAND2_X1 U789 ( .A1(G8), .A2(n690), .ZN(n691) );
  XNOR2_X1 U790 ( .A(KEYINPUT30), .B(n691), .ZN(n692) );
  NOR2_X1 U791 ( .A1(G168), .A2(n692), .ZN(n693) );
  NOR2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n696) );
  INV_X1 U793 ( .A(G1996), .ZN(n947) );
  XNOR2_X1 U794 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n697) );
  XNOR2_X1 U795 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n731), .A2(G1341), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U798 ( .A1(n701), .A2(n989), .ZN(n703) );
  OR2_X1 U799 ( .A1(n710), .A2(n977), .ZN(n709) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n714), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n704), .B(KEYINPUT96), .ZN(n706) );
  NAND2_X1 U802 ( .A1(G1348), .A2(n731), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U804 ( .A(KEYINPUT97), .B(n707), .Z(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n710), .A2(n977), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n714), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U809 ( .A(n713), .B(KEYINPUT27), .ZN(n716) );
  INV_X1 U810 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U811 ( .A1(n999), .A2(n714), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n971), .A2(n719), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U815 ( .A1(n971), .A2(n719), .ZN(n720) );
  XOR2_X1 U816 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(n723), .B(KEYINPUT29), .ZN(n726) );
  NOR2_X1 U819 ( .A1(G301), .A2(n724), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(KEYINPUT99), .ZN(n743) );
  AND2_X1 U823 ( .A1(G286), .A2(G8), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n743), .A2(n730), .ZN(n738) );
  INV_X1 U825 ( .A(G8), .ZN(n736) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n799), .ZN(n733) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n734), .A2(G303), .ZN(n735) );
  OR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  AND2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n740) );
  XOR2_X1 U832 ( .A(KEYINPUT32), .B(KEYINPUT100), .Z(n739) );
  NAND2_X1 U833 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n794) );
  NOR2_X1 U836 ( .A1(n796), .A2(n794), .ZN(n752) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n746) );
  XNOR2_X1 U838 ( .A(n746), .B(KEYINPUT101), .ZN(n748) );
  INV_X1 U839 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n750) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n793) );
  AND2_X1 U843 ( .A1(n981), .A2(KEYINPUT33), .ZN(n753) );
  INV_X1 U844 ( .A(n799), .ZN(n801) );
  NAND2_X1 U845 ( .A1(n753), .A2(n801), .ZN(n785) );
  NOR2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n823) );
  NAND2_X1 U847 ( .A1(n878), .A2(G104), .ZN(n756) );
  XNOR2_X1 U848 ( .A(n756), .B(KEYINPUT90), .ZN(n758) );
  NAND2_X1 U849 ( .A1(G140), .A2(n879), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U851 ( .A(KEYINPUT34), .B(n759), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G128), .A2(n882), .ZN(n761) );
  NAND2_X1 U853 ( .A1(G116), .A2(n883), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U855 ( .A(KEYINPUT35), .B(n762), .Z(n763) );
  NOR2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U857 ( .A(KEYINPUT36), .B(n765), .ZN(n864) );
  XNOR2_X1 U858 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U859 ( .A1(n864), .A2(n814), .ZN(n931) );
  NAND2_X1 U860 ( .A1(n823), .A2(n931), .ZN(n820) );
  NAND2_X1 U861 ( .A1(n878), .A2(G105), .ZN(n767) );
  XNOR2_X1 U862 ( .A(KEYINPUT38), .B(KEYINPUT92), .ZN(n766) );
  XNOR2_X1 U863 ( .A(n767), .B(n766), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G141), .A2(n879), .ZN(n769) );
  NAND2_X1 U865 ( .A1(G129), .A2(n882), .ZN(n768) );
  NAND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U867 ( .A1(G117), .A2(n883), .ZN(n770) );
  XNOR2_X1 U868 ( .A(KEYINPUT91), .B(n770), .ZN(n771) );
  NOR2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n889) );
  AND2_X1 U871 ( .A1(n889), .A2(G1996), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G95), .A2(n878), .ZN(n776) );
  NAND2_X1 U873 ( .A1(G131), .A2(n879), .ZN(n775) );
  NAND2_X1 U874 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G119), .A2(n882), .ZN(n778) );
  NAND2_X1 U876 ( .A1(G107), .A2(n883), .ZN(n777) );
  NAND2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n874) );
  INV_X1 U879 ( .A(G1991), .ZN(n955) );
  NOR2_X1 U880 ( .A1(n874), .A2(n955), .ZN(n781) );
  NOR2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n921) );
  INV_X1 U882 ( .A(n823), .ZN(n783) );
  NOR2_X1 U883 ( .A1(n921), .A2(n783), .ZN(n817) );
  INV_X1 U884 ( .A(n817), .ZN(n784) );
  AND2_X1 U885 ( .A1(n820), .A2(n784), .ZN(n808) );
  NAND2_X1 U886 ( .A1(n785), .A2(n808), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G1976), .A2(G288), .ZN(n979) );
  INV_X1 U888 ( .A(n979), .ZN(n786) );
  NOR2_X1 U889 ( .A1(n799), .A2(n786), .ZN(n787) );
  OR2_X1 U890 ( .A1(KEYINPUT33), .A2(n787), .ZN(n789) );
  XNOR2_X1 U891 ( .A(G1981), .B(G305), .ZN(n991) );
  INV_X1 U892 ( .A(n991), .ZN(n788) );
  NAND2_X1 U893 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U894 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U895 ( .A1(n793), .A2(n792), .ZN(n810) );
  OR2_X1 U896 ( .A1(n794), .A2(n801), .ZN(n795) );
  NAND2_X1 U897 ( .A1(G166), .A2(G8), .ZN(n797) );
  NOR2_X1 U898 ( .A1(G2090), .A2(n797), .ZN(n798) );
  AND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n804) );
  NOR2_X1 U900 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XNOR2_X1 U901 ( .A(n800), .B(KEYINPUT24), .ZN(n802) );
  AND2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X2 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT102), .ZN(n813) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n974) );
  NAND2_X1 U909 ( .A1(n974), .A2(n823), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n826) );
  NAND2_X1 U911 ( .A1(n864), .A2(n814), .ZN(n928) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n889), .ZN(n925) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n815) );
  AND2_X1 U914 ( .A1(n955), .A2(n874), .ZN(n923) );
  NOR2_X1 U915 ( .A1(n815), .A2(n923), .ZN(n816) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U917 ( .A1(n925), .A2(n818), .ZN(n819) );
  XNOR2_X1 U918 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n928), .A2(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G188) );
  XOR2_X1 U929 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n834), .ZN(G319) );
  XOR2_X1 U936 ( .A(KEYINPUT42), .B(G2078), .Z(n836) );
  XNOR2_X1 U937 ( .A(G2090), .B(G2084), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n837), .B(G2100), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U942 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U943 ( .A(KEYINPUT105), .B(G2678), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U945 ( .A(n843), .B(n842), .Z(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1966), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n846), .B(KEYINPUT107), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1971), .B(G1976), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1981), .B(G1956), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT106), .B(G2474), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G124), .A2(n882), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n855), .B(KEYINPUT44), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n856), .B(KEYINPUT108), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G100), .A2(n878), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G136), .A2(n879), .ZN(n860) );
  NAND2_X1 U964 ( .A1(G112), .A2(n883), .ZN(n859) );
  NAND2_X1 U965 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U966 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U967 ( .A(G164), .B(G160), .Z(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n895) );
  NAND2_X1 U969 ( .A1(n879), .A2(G142), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n865), .B(KEYINPUT110), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G106), .A2(n878), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT45), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G118), .A2(n883), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G130), .A2(n882), .ZN(n871) );
  XNOR2_X1 U977 ( .A(KEYINPUT109), .B(n871), .ZN(n872) );
  NOR2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n893) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n876) );
  XNOR2_X1 U980 ( .A(n874), .B(n919), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U982 ( .A(n877), .B(G162), .Z(n891) );
  NAND2_X1 U983 ( .A1(G103), .A2(n878), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G139), .A2(n879), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n882), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n934) );
  XOR2_X1 U991 ( .A(n889), .B(n934), .Z(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(n893), .B(n892), .Z(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U995 ( .A1(G37), .A2(n896), .ZN(G395) );
  INV_X1 U996 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U997 ( .A(G171), .B(n977), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(G286), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2454), .B(G2435), .Z(n902) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2427), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n902), .B(n901), .ZN(n909) );
  XOR2_X1 U1004 ( .A(KEYINPUT103), .B(G2446), .Z(n904) );
  XNOR2_X1 U1005 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U1006 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1007 ( .A(n905), .B(G2451), .Z(n907) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n910), .A2(G14), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(G2084), .B(G160), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(KEYINPUT111), .B(n917), .ZN(n918) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT112), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n939) );
  XOR2_X1 U1032 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n937), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n940), .ZN(n942) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n943), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1041 ( .A(G29), .B(KEYINPUT118), .Z(n969) );
  XNOR2_X1 U1042 ( .A(G2084), .B(G34), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(KEYINPUT54), .ZN(n966) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G32), .B(n947), .ZN(n948) );
  NAND2_X1 U1048 ( .A1(n948), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G27), .B(n949), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(KEYINPUT114), .B(n950), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1053 ( .A(n955), .B(G25), .Z(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1055 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT116), .B(n958), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n960), .B(n959), .ZN(n963) );
  XOR2_X1 U1058 ( .A(G2090), .B(G35), .Z(n961) );
  XNOR2_X1 U1059 ( .A(KEYINPUT113), .B(n961), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n964), .B(KEYINPUT117), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(n967), .B(KEYINPUT55), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n970), .ZN(n1030) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1067 ( .A(G171), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT120), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(n972), .B(n999), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(G1348), .B(KEYINPUT119), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(n977), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G166), .B(G1971), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1077 ( .A(KEYINPUT121), .B(n983), .Z(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n988), .ZN(n996) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1341), .ZN(n994) );
  XOR2_X1 U1082 ( .A(G1966), .B(G168), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT57), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1028) );
  INV_X1 U1088 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1089 ( .A(G20), .B(n999), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT123), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G6), .B(G1981), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(G4), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT60), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(KEYINPUT125), .B(n1010), .Z(n1012) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1013), .ZN(n1023) );
  XNOR2_X1 U1104 ( .A(n1014), .B(G5), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1110 ( .A(n1019), .B(KEYINPUT58), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(n1033), .B(KEYINPUT62), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1034), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

