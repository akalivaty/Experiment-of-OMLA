//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT83), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT66), .B1(new_n192), .B2(new_n194), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT5), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n192), .B2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n195), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G101), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n206), .B2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n206), .A3(G104), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(KEYINPUT80), .A3(G107), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n212), .A2(new_n214), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n211), .B1(new_n218), .B2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT82), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(new_n211), .C1(new_n218), .C2(G101), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT2), .B(G113), .Z(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n196), .B2(new_n200), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n199), .B1(new_n197), .B2(new_n198), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n190), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n192), .A2(new_n194), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n224), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n214), .A2(new_n217), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n212), .A4(new_n216), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n218), .A2(G101), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n218), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n223), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n223), .B(new_n244), .C1(new_n234), .C2(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT64), .B1(new_n251), .B2(G146), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(G143), .B2(new_n254), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n251), .A2(KEYINPUT65), .A3(G146), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n256), .B(new_n262), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n257), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(new_n251), .B2(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n254), .A3(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(KEYINPUT0), .A3(G128), .A4(new_n256), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G224), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n248), .A2(new_n250), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n244), .B(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n195), .B1(new_n204), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n220), .A2(new_n222), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n219), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n205), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n283), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT7), .B1(new_n279), .B2(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n278), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n290), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n269), .B(new_n292), .C1(new_n277), .C2(new_n268), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n247), .A2(new_n289), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT84), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n282), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n296), .A3(new_n299), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n298), .A2(KEYINPUT85), .A3(new_n300), .A4(new_n302), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT75), .A2(G125), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G140), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT76), .B1(new_n312), .B2(G125), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT75), .A3(G125), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT16), .A4(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n268), .A2(G140), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n315), .A2(KEYINPUT77), .ZN(new_n321));
  OAI21_X1  g135(.A(G146), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n313), .A2(new_n314), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n316), .A3(KEYINPUT16), .A4(new_n311), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n254), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(G237), .A2(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(G143), .A3(G214), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G143), .B1(new_n327), .B2(G214), .ZN(new_n330));
  OAI21_X1  g144(.A(G131), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n322), .A2(KEYINPUT87), .A3(new_n333), .A4(new_n326), .ZN(new_n337));
  INV_X1    g151(.A(new_n330), .ZN(new_n338));
  INV_X1    g152(.A(G131), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n328), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n340), .A3(new_n332), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n337), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(G113), .B(G122), .Z(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT86), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n208), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n329), .A2(new_n330), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT18), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(new_n339), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n323), .A2(new_n311), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G146), .ZN(new_n353));
  INV_X1    g167(.A(new_n317), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n268), .A2(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n254), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n344), .A2(new_n347), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n347), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n331), .A2(new_n340), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n254), .B1(new_n324), .B2(new_n325), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT19), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n354), .A2(new_n363), .A3(new_n355), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n352), .B2(KEYINPUT19), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n361), .B(new_n362), .C1(new_n365), .C2(new_n254), .ZN(new_n366));
  INV_X1    g180(.A(new_n358), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G475), .B1(new_n359), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n369), .A2(KEYINPUT20), .A3(new_n295), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT20), .B1(new_n369), .B2(new_n295), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n344), .A2(new_n347), .A3(new_n358), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n347), .B1(new_n344), .B2(new_n358), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n295), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT89), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n295), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G475), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT90), .A2(G122), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT90), .A2(G122), .ZN(new_n382));
  OAI21_X1  g196(.A(G116), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n206), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n191), .A2(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G128), .B(G143), .ZN(new_n388));
  INV_X1    g202(.A(G134), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n386), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n261), .A2(KEYINPUT13), .A3(G143), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n393), .A2(new_n395), .B1(new_n389), .B2(new_n388), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n386), .A2(G107), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n206), .B1(new_n383), .B2(new_n385), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT9), .B(G234), .Z(new_n401));
  INV_X1    g215(.A(G953), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(G217), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n392), .A2(KEYINPUT91), .A3(new_n399), .A4(new_n406), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n295), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n380), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G234), .ZN(new_n415));
  INV_X1    g229(.A(G237), .ZN(new_n416));
  OAI211_X1 g230(.A(G902), .B(G953), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(KEYINPUT92), .Z(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT21), .B(G898), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n402), .A2(G952), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n415), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AND4_X1   g237(.A1(new_n189), .A2(new_n308), .A3(new_n414), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n260), .A2(new_n266), .A3(KEYINPUT69), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT69), .B1(new_n260), .B2(new_n266), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT10), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n220), .A2(new_n222), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT11), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n389), .B2(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n389), .A2(G137), .ZN(new_n433));
  INV_X1    g247(.A(G137), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n432), .A2(new_n435), .A3(new_n339), .A4(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT68), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(KEYINPUT68), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n266), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n275), .A2(new_n256), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n259), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n275), .A2(KEYINPUT81), .A3(new_n256), .A4(new_n262), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n287), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n239), .A2(new_n277), .A3(new_n241), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n430), .A2(new_n443), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n260), .A2(new_n266), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n220), .B2(new_n222), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n439), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT12), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G140), .ZN(new_n460));
  INV_X1    g274(.A(G227), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n460), .B(new_n462), .Z(new_n463));
  NOR2_X1   g277(.A1(new_n443), .A2(KEYINPUT12), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n455), .B2(new_n457), .ZN(new_n465));
  AND4_X1   g279(.A1(new_n454), .A2(new_n459), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n452), .A2(new_n453), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n428), .A2(new_n429), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n442), .B(new_n441), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n463), .B1(new_n469), .B2(new_n454), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n425), .B(new_n295), .C1(new_n466), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(G469), .A2(G902), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n454), .A2(new_n459), .A3(new_n465), .ZN(new_n473));
  INV_X1    g287(.A(new_n463), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n454), .A3(new_n463), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(G469), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n401), .ZN(new_n479));
  OAI21_X1  g293(.A(G221), .B1(new_n479), .B2(G902), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n193), .A2(G128), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n193), .B2(G128), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n261), .A2(KEYINPUT73), .A3(KEYINPUT23), .A4(G119), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G119), .B(G128), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT24), .B(G110), .Z(new_n491));
  OAI22_X1  g305(.A1(new_n489), .A2(G110), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n322), .A2(new_n356), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n490), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n324), .A2(new_n254), .A3(new_n325), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(new_n362), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n489), .A2(KEYINPUT74), .A3(G110), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT74), .B1(new_n489), .B2(G110), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n493), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n499), .B(new_n494), .C1(new_n495), .C2(new_n362), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT78), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n493), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n402), .A2(G221), .A3(G234), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT22), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G137), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n502), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n503), .A2(new_n504), .A3(new_n493), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n295), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  INV_X1    g328(.A(G217), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(G234), .B2(new_n295), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n517), .A3(new_n295), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT79), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n521), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n516), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n481), .A2(new_n520), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n433), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n389), .A2(G137), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n438), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n426), .B2(new_n427), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n441), .A2(new_n277), .A3(new_n442), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n234), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n277), .A2(new_n439), .B1(new_n456), .B2(new_n530), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n234), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n439), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n272), .A2(new_n276), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n267), .B2(new_n529), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT67), .B1(new_n225), .B2(new_n195), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n230), .A2(new_n227), .A3(new_n232), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT71), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n533), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n535), .B1(KEYINPUT28), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(G101), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n327), .A2(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n544), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n533), .ZN(new_n557));
  INV_X1    g371(.A(new_n551), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT72), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n552), .A2(new_n559), .A3(new_n562), .A4(new_n553), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n531), .A2(new_n532), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n544), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n533), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n535), .B1(KEYINPUT28), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n558), .A2(new_n553), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n533), .A2(new_n551), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n533), .A2(KEYINPUT70), .A3(new_n551), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n574), .A2(new_n556), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n547), .B2(new_n551), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n533), .A2(KEYINPUT70), .A3(new_n551), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT70), .B1(new_n533), .B2(new_n551), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n575), .B1(new_n581), .B2(new_n556), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n571), .B(new_n295), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT32), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n556), .A3(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT31), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n577), .C1(new_n551), .C2(new_n547), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n571), .A4(new_n295), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n570), .A2(G472), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n525), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n424), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NAND2_X1  g407(.A1(new_n583), .A2(KEYINPUT93), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n571), .B1(new_n587), .B2(new_n295), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT93), .B(new_n571), .C1(new_n587), .C2(new_n295), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n525), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n408), .A2(new_n409), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n404), .A2(KEYINPUT33), .A3(new_n407), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n411), .A2(G902), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n604), .A2(new_n605), .B1(new_n411), .B2(new_n410), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n380), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n423), .ZN(new_n609));
  INV_X1    g423(.A(new_n306), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n299), .B1(new_n282), .B2(new_n296), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n189), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n599), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n297), .A2(new_n300), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n188), .B1(new_n617), .B2(new_n306), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n618), .A2(new_n372), .A3(new_n413), .A4(new_n379), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n423), .B(KEYINPUT94), .Z(new_n620));
  OR3_X1    g434(.A1(new_n619), .A2(KEYINPUT95), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT95), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n623), .A2(new_n525), .A3(new_n598), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  INV_X1    g440(.A(new_n598), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n501), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n523), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n520), .A2(new_n522), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n481), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n424), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT37), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(G12));
  NAND2_X1  g449(.A1(new_n570), .A2(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n584), .A2(new_n589), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g452(.A1(new_n638), .A2(new_n481), .A3(new_n618), .A4(new_n631), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n372), .A2(new_n413), .A3(new_n379), .ZN(new_n640));
  INV_X1    g454(.A(new_n422), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n418), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XNOR2_X1  g461(.A(new_n643), .B(KEYINPUT98), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT39), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n481), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n581), .A2(new_n556), .B1(new_n558), .B2(new_n566), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n653), .B2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT96), .ZN(new_n656));
  INV_X1    g470(.A(new_n631), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n308), .B(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n380), .A2(new_n413), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n188), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n651), .B(new_n652), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT99), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n661), .B(KEYINPUT97), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n651), .A4(new_n652), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n251), .ZN(G45));
  AOI211_X1 g484(.A(new_n643), .B(new_n606), .C1(new_n372), .C2(new_n379), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n639), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AND3_X1   g487(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n295), .B1(new_n466), .B2(new_n470), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n480), .A3(new_n471), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n613), .A2(new_n638), .A3(new_n674), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND3_X1  g495(.A1(new_n674), .A2(new_n638), .A3(new_n678), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n623), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n191), .ZN(G18));
  AND2_X1   g498(.A1(new_n631), .A2(new_n414), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n677), .A2(new_n612), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n423), .A3(new_n638), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NOR3_X1   g502(.A1(new_n659), .A2(new_n612), .A3(new_n677), .ZN(new_n689));
  INV_X1    g503(.A(new_n620), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n577), .B1(new_n567), .B2(new_n551), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n571), .B(new_n295), .C1(new_n691), .C2(new_n582), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n595), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n674), .A3(new_n690), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NAND4_X1  g510(.A1(new_n631), .A2(new_n671), .A3(new_n694), .A4(new_n686), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  AND4_X1   g516(.A1(new_n189), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n475), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n473), .A2(KEYINPUT102), .A3(new_n474), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(G469), .A3(new_n476), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n472), .B(KEYINPUT101), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n471), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n480), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n703), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n305), .A2(new_n189), .A3(new_n306), .A4(new_n307), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT103), .B1(new_n714), .B2(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n674), .A2(new_n638), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n671), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n671), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n722), .B(new_n717), .C1(new_n713), .C2(new_n715), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n721), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NAND3_X1  g541(.A1(new_n716), .A2(new_n645), .A3(new_n718), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  INV_X1    g543(.A(new_n380), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n607), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(KEYINPUT43), .Z(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n598), .A3(new_n631), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n475), .B2(new_n476), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n425), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n476), .A4(new_n707), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n709), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(KEYINPUT105), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n471), .ZN(new_n743));
  INV_X1    g557(.A(new_n709), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n737), .B2(new_n738), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n743), .B1(new_n745), .B2(KEYINPUT46), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n745), .B2(KEYINPUT46), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n742), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n480), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n649), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n714), .B1(new_n733), .B2(new_n734), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n735), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n434), .ZN(G39));
  AND3_X1   g569(.A1(new_n749), .A2(KEYINPUT106), .A3(new_n480), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT106), .B1(new_n749), .B2(new_n480), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  OAI22_X1  g577(.A1(new_n756), .A2(new_n760), .B1(new_n763), .B2(KEYINPUT47), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n762), .A2(new_n764), .A3(new_n703), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n674), .A2(new_n638), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n671), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n764), .A3(new_n671), .A4(new_n703), .ZN(new_n769));
  INV_X1    g583(.A(new_n767), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT108), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AND4_X1   g587(.A1(new_n641), .A2(new_n732), .A3(new_n674), .A4(new_n694), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n658), .A2(new_n189), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n678), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT50), .Z(new_n777));
  AND2_X1   g591(.A1(new_n762), .A2(new_n764), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n676), .A2(new_n471), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n480), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n703), .B(new_n774), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n674), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n656), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n714), .A2(new_n422), .A3(new_n677), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n730), .A3(new_n606), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n631), .A2(new_n694), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n732), .A2(new_n787), .A3(new_n785), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT114), .Z(new_n789));
  NAND4_X1  g603(.A1(new_n777), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT51), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n640), .A2(KEYINPUT110), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n380), .B2(new_n607), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n796), .B2(new_n640), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n308), .A2(new_n189), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n599), .A2(new_n797), .A3(new_n798), .A4(new_n690), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n633), .A3(new_n687), .A4(new_n592), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n679), .B(new_n695), .C1(new_n623), .C2(new_n682), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n726), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  INV_X1    g618(.A(new_n608), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n704), .B1(new_n703), .B2(new_n712), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n714), .A2(KEYINPUT103), .A3(new_n711), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n805), .B(new_n787), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n638), .A2(new_n481), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n631), .A2(new_n414), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n714), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n643), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n728), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n804), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n608), .B1(new_n713), .B2(new_n715), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n811), .B1(new_n816), .B2(new_n787), .ZN(new_n817));
  OAI211_X1 g631(.A(KEYINPUT111), .B(new_n728), .C1(new_n817), .C2(new_n643), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n803), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n699), .A2(new_n700), .B1(new_n645), .B2(new_n639), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n520), .A2(new_n522), .A3(new_n630), .A4(new_n644), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT112), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n610), .A2(new_n611), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n659), .A2(new_n188), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n656), .A3(new_n712), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(new_n700), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n672), .B(new_n646), .C1(new_n828), .C2(new_n698), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n821), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n655), .A2(KEYINPUT96), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT96), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n637), .B2(new_n654), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n824), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n831), .A2(new_n835), .A3(new_n711), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n827), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n819), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n815), .A2(new_n818), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n802), .A2(new_n726), .ZN(new_n841));
  AND4_X1   g655(.A1(KEYINPUT53), .A2(new_n840), .A3(new_n841), .A4(new_n838), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n793), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n838), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n841), .A3(new_n838), .A4(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n784), .A2(new_n805), .A3(new_n785), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n732), .A2(new_n718), .A3(new_n785), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  AOI211_X1 g666(.A(new_n850), .B(new_n852), .C1(new_n686), .C2(new_n774), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n421), .A3(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n792), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n658), .A2(new_n188), .A3(new_n731), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n779), .B(KEYINPUT49), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n784), .A3(new_n480), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT109), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(G75));
  AOI21_X1  g674(.A(new_n295), .B1(new_n846), .B2(new_n847), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(G210), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n248), .A2(new_n250), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(new_n281), .Z(new_n866));
  XOR2_X1   g680(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n864), .A2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n402), .A2(G952), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G51));
  XOR2_X1   g687(.A(new_n709), .B(KEYINPUT57), .Z(new_n874));
  NAND3_X1  g688(.A1(new_n843), .A2(new_n848), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n843), .A2(new_n877), .A3(new_n848), .A4(new_n874), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n876), .B(new_n878), .C1(new_n470), .C2(new_n466), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n861), .A2(new_n738), .A3(new_n737), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n872), .B1(new_n879), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n861), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n359), .A2(new_n368), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n882), .A2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n872), .ZN(G60));
  XNOR2_X1  g701(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n411), .A2(new_n295), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n843), .A2(new_n848), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(new_n603), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n603), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n872), .ZN(G63));
  XNOR2_X1  g708(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n515), .A2(new_n295), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n629), .B(new_n897), .C1(new_n839), .C2(new_n842), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n901));
  INV_X1    g715(.A(new_n897), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n846), .B2(new_n847), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n629), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n872), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n903), .B2(new_n512), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n906), .C1(new_n903), .C2(new_n512), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n900), .A2(new_n904), .B1(new_n901), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(G66));
  OAI21_X1  g731(.A(G953), .B1(new_n419), .B2(new_n279), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n802), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n865), .B1(G898), .B2(new_n402), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  OAI21_X1  g735(.A(G953), .B1(new_n461), .B2(new_n642), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT125), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n554), .A2(new_n555), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n365), .B(KEYINPUT123), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  INV_X1    g742(.A(new_n829), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n665), .A2(new_n668), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n665), .A2(new_n668), .A3(KEYINPUT62), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n754), .B1(new_n768), .B2(new_n771), .ZN(new_n935));
  INV_X1    g749(.A(new_n797), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n936), .A2(new_n717), .A3(new_n650), .A4(new_n714), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n928), .B1(new_n939), .B2(new_n402), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n752), .A2(new_n718), .A3(new_n824), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n726), .A2(new_n929), .A3(new_n728), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n935), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n402), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n402), .A2(G900), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n927), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n924), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n927), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n941), .B(new_n754), .C1(new_n768), .C2(new_n771), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n951), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n946), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n937), .B1(new_n932), .B2(new_n933), .ZN(new_n954));
  AOI21_X1  g768(.A(G953), .B1(new_n954), .B2(new_n935), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n953), .B(new_n923), .C1(new_n955), .C2(new_n928), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n949), .A2(new_n956), .ZN(G72));
  XNOR2_X1  g771(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n958));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n802), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n944), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n557), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n558), .A3(new_n963), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n846), .A2(new_n847), .B1(new_n585), .B2(new_n559), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n872), .B1(new_n965), .B2(new_n960), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n934), .A2(new_n802), .A3(new_n935), .A4(new_n938), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n960), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n963), .A2(new_n558), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(KEYINPUT127), .A3(new_n970), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(G57));
endmodule


