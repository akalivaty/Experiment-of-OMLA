//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(new_n206), .B2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G13), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n219), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n216), .B(new_n223), .C1(new_n226), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n251), .A2(new_n252), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(G226), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT70), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n268), .B1(new_n208), .B2(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n224), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT71), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n225), .A2(KEYINPUT71), .A3(G33), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g0084(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n225), .A2(new_n279), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n285), .A2(new_n225), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n277), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n277), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n260), .A2(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G50), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n289), .B(new_n294), .C1(G50), .C2(new_n290), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n275), .B(new_n296), .C1(new_n297), .C2(new_n274), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n275), .B2(KEYINPUT74), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n298), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n274), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT72), .B(G179), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n265), .A2(new_n304), .A3(new_n273), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n291), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n292), .A2(G68), .A3(new_n293), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n282), .A2(new_n208), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G50), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n225), .B2(G68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(KEYINPUT75), .B2(new_n314), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n277), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT11), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n310), .B(new_n311), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n266), .A2(G226), .A3(new_n267), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n269), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n272), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n258), .B1(G238), .B2(new_n263), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n325), .B(G169), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G179), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n325), .B1(new_n341), .B2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n324), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G200), .B1(new_n333), .B2(new_n334), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(G190), .A3(new_n338), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n323), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n283), .B1(new_n260), .B2(G20), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n292), .B1(new_n291), .B2(new_n283), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n277), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G33), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT7), .B1(new_n356), .B2(new_n225), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n358), .B(G20), .C1(new_n353), .C2(new_n355), .ZN(new_n359));
  OAI21_X1  g0159(.A(G68), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G58), .A2(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n227), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n313), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n352), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(KEYINPUT77), .A3(new_n364), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT77), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n225), .B1(new_n227), .B2(new_n361), .ZN(new_n372));
  INV_X1    g0172(.A(new_n364), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT16), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n356), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n266), .A2(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n225), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n359), .B1(new_n379), .B2(new_n358), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n380), .B2(new_n308), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n351), .B1(new_n369), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n259), .A2(G232), .A3(new_n261), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n257), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n353), .A2(new_n355), .A3(G223), .A4(new_n267), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n353), .A2(new_n355), .A3(G226), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n272), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n304), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n272), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n257), .A2(new_n383), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G169), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT18), .B1(new_n382), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n393), .A3(new_n297), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n389), .B2(G200), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT16), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT76), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT76), .B1(new_n353), .B2(new_n355), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(G20), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(KEYINPUT7), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n406), .B2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n358), .B1(new_n266), .B2(G20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n402), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n365), .B1(new_n409), .B2(G68), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n277), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n350), .B(new_n400), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n350), .B1(new_n407), .B2(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(new_n396), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n369), .A2(new_n381), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n350), .A4(new_n400), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n398), .A2(new_n414), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT15), .B(G87), .Z(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n282), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n283), .A2(new_n286), .B1(new_n225), .B2(new_n208), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n277), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n352), .A2(new_n290), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n293), .A2(G77), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT73), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n292), .A2(new_n429), .A3(G77), .A4(new_n293), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n425), .B(new_n431), .C1(G77), .C2(new_n290), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n257), .B1(new_n262), .B2(new_n207), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n434));
  INV_X1    g0234(.A(G238), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n203), .B2(new_n266), .C1(new_n269), .C2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n436), .B2(new_n272), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(G190), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n437), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n437), .A2(G169), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n304), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n432), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n307), .A2(new_n348), .A3(new_n420), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n260), .A2(G33), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n290), .A2(new_n446), .A3(new_n224), .A4(new_n276), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT25), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n290), .B2(G107), .ZN(new_n451));
  AOI22_X1  g0251(.A1(G107), .A2(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT23), .B1(new_n203), .B2(G20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n454), .A2(new_n455), .B1(G20), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n353), .A2(new_n355), .A3(new_n225), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n266), .A2(new_n460), .A3(new_n225), .A4(G87), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n453), .B1(new_n464), .B2(new_n277), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  INV_X1    g0266(.A(G294), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n279), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G250), .A2(G1698), .ZN(new_n469));
  INV_X1    g0269(.A(G257), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(G1698), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n266), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n466), .B1(new_n472), .B2(new_n259), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n255), .A2(G1), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G264), .A3(new_n259), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n253), .A2(new_n479), .A3(new_n474), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n468), .ZN(new_n482));
  OR2_X1    g0282(.A1(G250), .A2(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(G1698), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n356), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT84), .A3(new_n272), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n473), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n272), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n489), .A2(new_n478), .A3(new_n480), .ZN(new_n490));
  AOI22_X1  g0290(.A1(G169), .A2(new_n488), .B1(new_n490), .B2(G179), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT85), .B1(new_n465), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(KEYINPUT24), .B(new_n457), .C1(new_n459), .C2(new_n461), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n459), .A2(new_n461), .ZN(new_n494));
  INV_X1    g0294(.A(new_n457), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n463), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n277), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n452), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(G169), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n490), .A2(G179), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n447), .A2(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n291), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n276), .A2(new_n224), .B1(G20), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n225), .C1(G33), .C2(new_n202), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n509), .A2(KEYINPUT20), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT20), .B1(new_n509), .B2(new_n511), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n506), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G169), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n477), .A2(G270), .A3(new_n259), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n480), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n353), .A2(new_n355), .A3(G264), .A4(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n266), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n356), .A2(G303), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n266), .A2(G257), .A3(new_n267), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n517), .B1(new_n524), .B2(new_n272), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n515), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n525), .A2(G179), .A3(new_n514), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n505), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n272), .ZN(new_n530));
  INV_X1    g0330(.A(new_n517), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(KEYINPUT21), .A3(G169), .A4(new_n514), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n525), .A2(G179), .A3(new_n514), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(KEYINPUT83), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n526), .B1(new_n515), .B2(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n504), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n272), .B1(new_n474), .B2(new_n479), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n272), .A2(new_n486), .B1(new_n539), .B2(G264), .ZN(new_n540));
  AOI21_X1  g0340(.A(G200), .B1(new_n540), .B2(new_n480), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n297), .A2(new_n473), .A3(new_n481), .A4(new_n487), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(KEYINPUT86), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n488), .B2(G190), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n498), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n548), .A2(new_n202), .A3(G107), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n313), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n409), .A2(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n352), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n290), .A2(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n448), .B2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n477), .A2(G257), .A3(new_n259), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n480), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n353), .A2(new_n355), .A3(G244), .A4(new_n267), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n510), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n566), .B2(new_n272), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n555), .A2(new_n558), .B1(new_n567), .B2(G169), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n304), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n550), .B1(new_n547), .B2(new_n548), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(new_n225), .B1(new_n208), .B2(new_n286), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n203), .B1(new_n408), .B2(new_n402), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n277), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n557), .C1(new_n567), .C2(new_n439), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n567), .A2(G190), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n568), .A2(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n546), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n435), .A2(new_n267), .ZN(new_n579));
  INV_X1    g0379(.A(G244), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n353), .A2(new_n579), .A3(new_n355), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n456), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(KEYINPUT79), .A3(new_n456), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n259), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT78), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n253), .A2(new_n588), .A3(new_n474), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n253), .B2(new_n474), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n260), .A2(G45), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G250), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n590), .A2(new_n591), .B1(new_n272), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n587), .A2(new_n594), .A3(KEYINPUT80), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT80), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n582), .A2(KEYINPUT79), .A3(new_n456), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT79), .B1(new_n582), .B2(new_n456), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n272), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n272), .A2(new_n593), .ZN(new_n600));
  INV_X1    g0400(.A(new_n591), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n589), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n302), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT80), .B1(new_n587), .B2(new_n594), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n602), .A3(new_n596), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n304), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n421), .A2(new_n290), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n266), .A2(new_n225), .A3(G68), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n225), .B1(new_n327), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(G87), .B2(new_n204), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n202), .B1(new_n280), .B2(new_n281), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n609), .B(new_n612), .C1(new_n613), .C2(KEYINPUT19), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n352), .B1(new_n614), .B2(KEYINPUT81), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n610), .B1(new_n282), .B2(new_n202), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT81), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n609), .A4(new_n612), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n608), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n448), .A2(new_n421), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n604), .A2(new_n607), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(G200), .B1(new_n595), .B2(new_n603), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n605), .A2(G190), .A3(new_n606), .ZN(new_n624));
  INV_X1    g0424(.A(G87), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n447), .A2(new_n625), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n608), .B(new_n626), .C1(new_n615), .C2(new_n618), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n514), .B1(new_n525), .B2(G190), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n439), .B2(new_n525), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n622), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n445), .A2(new_n538), .A3(new_n578), .A4(new_n631), .ZN(G372));
  OAI21_X1  g0432(.A(new_n302), .B1(new_n587), .B2(new_n594), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n607), .A2(new_n621), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(G200), .B1(new_n587), .B2(new_n594), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n624), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n568), .A2(new_n570), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n622), .A2(new_n628), .A3(KEYINPUT26), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n634), .A2(new_n636), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n527), .A2(new_n528), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n498), .A2(new_n501), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .A4(new_n536), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n533), .A2(new_n536), .A3(new_n534), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n497), .A2(new_n452), .B1(new_n499), .B2(new_n500), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT87), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n643), .A2(new_n578), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n651), .A3(new_n634), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n445), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n306), .ZN(new_n654));
  INV_X1    g0454(.A(new_n443), .ZN(new_n655));
  OAI21_X1  g0455(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n339), .A3(new_n335), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n324), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n347), .A2(new_n414), .A3(new_n419), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n398), .B(new_n417), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n661), .B2(new_n301), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n653), .A2(new_n662), .ZN(G369));
  NOR2_X1   g0463(.A1(new_n504), .A2(new_n546), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n260), .A2(new_n225), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(G213), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n664), .B1(new_n465), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n649), .A2(new_n670), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n514), .A2(new_n670), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n630), .B1(new_n648), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n537), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n537), .A2(new_n671), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(new_n664), .B1(new_n649), .B2(new_n671), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n221), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n229), .B2(new_n686), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n605), .A2(new_n540), .A3(new_n606), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n605), .A2(new_n695), .A3(new_n606), .A4(new_n540), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n566), .A2(new_n272), .ZN(new_n697));
  INV_X1    g0497(.A(new_n560), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G179), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n532), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n587), .B2(new_n594), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT89), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n705), .A2(new_n699), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n490), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n304), .A3(new_n532), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n703), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n702), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(new_n699), .A3(new_n706), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT30), .B1(new_n713), .B2(new_n709), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n694), .A3(new_n696), .A4(new_n701), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n671), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n670), .A3(new_n715), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n716), .A2(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n538), .A2(new_n631), .A3(new_n578), .A4(new_n671), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n692), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n652), .A2(new_n671), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT90), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n652), .A2(new_n726), .A3(new_n671), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n622), .A2(new_n628), .A3(new_n637), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT91), .A3(new_n639), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n637), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT91), .B1(new_n729), .B2(new_n639), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n634), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT92), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n538), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n737));
  INV_X1    g0537(.A(new_n541), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n545), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n465), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n634), .A3(new_n636), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n699), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n567), .A2(G190), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n574), .A3(new_n557), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n574), .A2(new_n557), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n569), .C1(G169), .C2(new_n567), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n743), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n741), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT92), .B1(new_n504), .B2(new_n537), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n736), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(KEYINPUT29), .B(new_n671), .C1(new_n734), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n722), .B1(new_n728), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n691), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n219), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n260), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n686), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n221), .A2(new_n266), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n221), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n248), .A2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n403), .A2(new_n404), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n221), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n255), .B2(new_n229), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n762), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n224), .B1(G20), .B2(new_n302), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n759), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n225), .A2(new_n297), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(new_n700), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n225), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G159), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n266), .B1(new_n625), .B2(new_n776), .C1(new_n781), .C2(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n390), .A2(G20), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n390), .A2(new_n439), .A3(new_n777), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n308), .B1(new_n208), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n782), .B(new_n787), .C1(KEYINPUT32), .C2(new_n781), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n777), .A2(new_n700), .A3(G200), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G107), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n783), .A2(new_n297), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n390), .A2(new_n439), .A3(new_n775), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n792), .A2(G50), .B1(new_n794), .B2(G58), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n225), .B1(new_n778), .B2(G190), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G97), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n788), .A2(new_n791), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n776), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n266), .B1(new_n800), .B2(G303), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n784), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n786), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G311), .A2(new_n805), .B1(new_n794), .B2(G322), .ZN(new_n806));
  INV_X1    g0606(.A(G329), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n807), .A2(new_n779), .B1(new_n796), .B2(new_n467), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n792), .B2(G326), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n790), .A2(G283), .B1(new_n801), .B2(KEYINPUT96), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n806), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n799), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n774), .B1(new_n812), .B2(new_n771), .ZN(new_n813));
  INV_X1    g0613(.A(new_n770), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n677), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n677), .A2(G330), .ZN(new_n816));
  INV_X1    g0616(.A(new_n759), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n678), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n443), .A2(KEYINPUT98), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n432), .A2(new_n670), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT98), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n441), .A2(new_n822), .A3(new_n442), .A4(new_n432), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n440), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n655), .A2(new_n670), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n724), .A2(new_n727), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n820), .A2(new_n440), .A3(new_n823), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n652), .A2(new_n671), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n722), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(KEYINPUT99), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(KEYINPUT99), .B2(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(new_n771), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n769), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n759), .B1(G77), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n356), .B1(new_n779), .B2(new_n838), .C1(new_n776), .C2(new_n203), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n790), .A2(G87), .ZN(new_n840));
  INV_X1    g0640(.A(new_n792), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n839), .B(new_n843), .C1(G294), .C2(new_n794), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n784), .A2(G283), .B1(new_n805), .B2(G116), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n798), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n794), .B1(new_n805), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n841), .B2(new_n849), .C1(new_n287), .C2(new_n785), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT34), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n790), .A2(G68), .ZN(new_n852));
  INV_X1    g0652(.A(new_n764), .ZN(new_n853));
  INV_X1    g0653(.A(new_n796), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G58), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n800), .A2(G50), .B1(new_n780), .B2(G132), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n847), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n837), .B1(new_n858), .B2(new_n771), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n824), .A2(new_n825), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n769), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n834), .A2(new_n861), .ZN(G384));
  XNOR2_X1  g0662(.A(new_n552), .B(KEYINPUT100), .ZN(new_n863));
  OAI211_X1 g0663(.A(G116), .B(new_n226), .C1(new_n863), .C2(KEYINPUT35), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(KEYINPUT101), .B1(KEYINPUT35), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT101), .B2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n361), .A2(G77), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n228), .A2(new_n868), .B1(G50), .B2(new_n308), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n219), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT102), .Z(new_n872));
  NAND3_X1  g0672(.A1(new_n728), .A2(new_n445), .A3(new_n753), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n662), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT105), .Z(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT7), .B1(new_n764), .B2(new_n225), .ZN(new_n877));
  OAI21_X1  g0677(.A(G68), .B1(new_n877), .B2(new_n359), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n352), .B1(new_n878), .B2(new_n375), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n379), .A2(new_n358), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n308), .B1(new_n880), .B2(new_n402), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n370), .A2(new_n374), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n368), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n351), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n668), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n412), .B1(new_n884), .B2(new_n397), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n886), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n415), .A2(new_n396), .ZN(new_n888));
  INV_X1    g0688(.A(new_n668), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n415), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n412), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n876), .B1(new_n420), .B2(new_n885), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n887), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n420), .A2(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n324), .A2(new_n670), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n343), .A2(new_n347), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n324), .B(new_n670), .C1(new_n658), .C2(new_n346), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n820), .A2(new_n823), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n671), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT103), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n829), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n398), .A2(new_n417), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n898), .A2(new_n907), .B1(new_n908), .B2(new_n668), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n412), .B1(new_n382), .B2(new_n397), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n382), .A2(new_n668), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n892), .A2(new_n913), .B1(new_n420), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n910), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n892), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n414), .A2(new_n419), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n912), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT104), .A3(new_n876), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n658), .A2(new_n324), .A3(new_n671), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n909), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n875), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n719), .A2(new_n717), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n721), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n826), .B1(new_n900), .B2(new_n901), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n893), .C2(new_n896), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n902), .A2(new_n860), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n720), .B2(new_n721), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n922), .A3(KEYINPUT40), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n445), .A2(new_n934), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n692), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n931), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n945), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n930), .A2(new_n947), .B1(new_n260), .B2(new_n756), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n872), .B1(new_n946), .B2(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n238), .A2(new_n765), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n772), .B1(new_n221), .B2(new_n422), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n759), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n797), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n308), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n792), .A2(G143), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n794), .A2(G150), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n789), .A2(new_n208), .B1(new_n779), .B2(new_n849), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n356), .B(new_n958), .C1(G58), .C2(new_n800), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n784), .A2(G159), .B1(new_n805), .B2(G50), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT108), .ZN(new_n962));
  INV_X1    g0762(.A(new_n789), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(G97), .B1(new_n780), .B2(G317), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n854), .A2(G107), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n800), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  AND4_X1   g0766(.A1(new_n764), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT46), .B1(new_n800), .B2(G116), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(KEYINPUT107), .B2(new_n968), .C1(new_n467), .C2(new_n785), .ZN(new_n969));
  AOI22_X1  g0769(.A1(KEYINPUT107), .A2(new_n968), .B1(new_n794), .B2(G303), .ZN(new_n970));
  INV_X1    g0770(.A(G283), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n970), .B1(new_n971), .B2(new_n786), .C1(new_n838), .C2(new_n841), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n960), .A2(new_n962), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n952), .B1(new_n974), .B2(new_n771), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n643), .B1(new_n627), .B2(new_n671), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n634), .A2(new_n627), .A3(new_n671), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n975), .B1(new_n978), .B2(new_n814), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n742), .A2(new_n749), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n747), .A2(new_n670), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n980), .A2(new_n981), .B1(new_n637), .B2(new_n670), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n683), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n983), .A2(new_n683), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n983), .B2(new_n683), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n680), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n986), .A2(new_n990), .A3(new_n680), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT106), .B1(new_n674), .B2(new_n682), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n682), .A2(new_n664), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n672), .A2(new_n998), .A3(new_n673), .A4(new_n681), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n679), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n678), .A3(new_n997), .A4(new_n999), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n754), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n754), .B1(new_n995), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n686), .B(KEYINPUT41), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n758), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n982), .A2(new_n997), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT42), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n980), .A2(new_n504), .A3(new_n981), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n670), .B1(new_n1010), .B2(new_n748), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n1008), .B2(KEYINPUT42), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n978), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1009), .A2(new_n1012), .A3(new_n1015), .A4(new_n1014), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n680), .A2(new_n982), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1020), .B(new_n1021), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n979), .B1(new_n1007), .B2(new_n1022), .ZN(G387));
  NAND3_X1  g0823(.A1(new_n672), .A2(new_n673), .A3(new_n770), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n234), .A2(new_n255), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1025), .A2(new_n765), .B1(new_n688), .B2(new_n760), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n688), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(new_n203), .B2(new_n685), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n759), .B1(new_n1031), .B2(new_n773), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n800), .A2(G77), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n853), .B(new_n1033), .C1(new_n287), .C2(new_n779), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G50), .B2(new_n794), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n792), .A2(G159), .B1(new_n805), .B2(G68), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n283), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n784), .B1(new_n790), .B2(G97), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n797), .A2(new_n421), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n963), .A2(G116), .B1(new_n780), .B2(G326), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n776), .A2(new_n467), .B1(new_n796), .B2(new_n971), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT109), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G303), .A2(new_n805), .B1(new_n794), .B2(G317), .ZN(new_n1044));
  INV_X1    g0844(.A(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n841), .B2(new_n1045), .C1(new_n838), .C2(new_n785), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n764), .B(new_n1041), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1040), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1032), .B1(new_n1053), .B2(new_n771), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1003), .A2(new_n758), .B1(new_n1024), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1004), .A2(new_n686), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1003), .A2(new_n754), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  AOI21_X1  g0858(.A(new_n757), .B1(new_n995), .B2(KEYINPUT110), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT110), .B2(new_n995), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n244), .A2(new_n765), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n772), .B1(new_n202), .B2(new_n221), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n759), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n792), .A2(G150), .B1(new_n794), .B2(G159), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT51), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n800), .A2(G68), .B1(new_n780), .B2(G143), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(new_n853), .A3(new_n840), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(G50), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n785), .A2(new_n1068), .B1(new_n283), .B2(new_n786), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n953), .A2(new_n208), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT111), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n792), .A2(G317), .B1(new_n794), .B2(G311), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n791), .B1(new_n467), .B2(new_n786), .C1(new_n785), .C2(new_n842), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n796), .A2(new_n508), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n356), .B1(new_n779), .B2(new_n1045), .C1(new_n776), .C2(new_n971), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1067), .A2(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n771), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n983), .B2(new_n814), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1060), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n995), .A2(new_n1004), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n995), .A2(new_n1004), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n686), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(new_n1085), .ZN(G390));
  NAND4_X1  g0886(.A1(new_n934), .A2(G330), .A3(new_n860), .A4(new_n902), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n922), .A2(new_n926), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n671), .B(new_n828), .C1(new_n734), .C2(new_n752), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n905), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n1091), .B2(new_n902), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n829), .A2(new_n906), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n902), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n926), .A2(new_n1094), .B1(new_n924), .B2(new_n925), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1088), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT38), .B1(new_n916), .B2(new_n918), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n887), .A2(new_n892), .B1(new_n420), .B2(new_n885), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(KEYINPUT104), .A2(new_n1097), .B1(new_n1098), .B2(KEYINPUT38), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n915), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n893), .A2(new_n896), .A3(new_n923), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n907), .B2(new_n927), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n903), .B1(new_n1090), .B2(new_n905), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1087), .C1(new_n1103), .C2(new_n1089), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1096), .A2(new_n758), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G97), .A2(new_n805), .B1(new_n794), .B2(G116), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n841), .B2(new_n971), .C1(new_n203), .C2(new_n785), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n852), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n356), .B1(new_n779), .B2(new_n467), .C1(new_n776), .C2(new_n625), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1070), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n780), .A2(G125), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n356), .B1(new_n963), .B2(G50), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1112), .C1(new_n841), .C2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n776), .A2(new_n287), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT114), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1114), .B(new_n1117), .C1(G132), .C2(new_n794), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n784), .A2(G137), .B1(new_n805), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(G159), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n953), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT113), .Z(new_n1124));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n759), .B1(new_n1037), .B2(new_n836), .C1(new_n1125), .C2(new_n835), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n924), .A2(new_n925), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n768), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1105), .A2(new_n1130), .A3(KEYINPUT116), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT116), .B1(new_n1105), .B2(new_n1130), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n829), .A2(new_n906), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n934), .A2(G330), .A3(new_n860), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n903), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1136), .B2(new_n1087), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1091), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1136), .A2(new_n1087), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n445), .A2(new_n722), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n873), .A2(new_n662), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT112), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n873), .A2(new_n662), .A3(new_n1141), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1136), .A2(new_n1087), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1093), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1136), .A2(new_n1090), .A3(new_n905), .A4(new_n1087), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT112), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1133), .A2(new_n1143), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1096), .A2(new_n1104), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n686), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1131), .A2(new_n1132), .B1(new_n1152), .B2(new_n1154), .ZN(G378));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1144), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n938), .A2(new_n941), .A3(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT118), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n692), .B1(new_n936), .B2(new_n937), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n941), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n295), .A2(new_n889), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n301), .A2(new_n306), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n301), .B2(new_n306), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1158), .A2(new_n1161), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n929), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1157), .A2(KEYINPUT118), .A3(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1161), .A2(new_n1172), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1160), .B1(new_n1159), .B2(new_n941), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1175), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n929), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1156), .A2(KEYINPUT57), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n686), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1174), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1156), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1181), .A2(new_n758), .A3(new_n1176), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n759), .B1(G50), .B2(new_n836), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n841), .A2(new_n508), .B1(new_n422), .B2(new_n786), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n784), .A2(G97), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n963), .A2(G58), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n780), .A2(G283), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(new_n1033), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n853), .A2(G41), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n203), .B2(new_n793), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1191), .A2(new_n1195), .A3(new_n1197), .A4(new_n954), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT58), .Z(new_n1199));
  OAI21_X1  g0999(.A(new_n1068), .B1(G33), .B2(G41), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1113), .A2(new_n793), .B1(new_n786), .B2(new_n849), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n784), .A2(G132), .B1(new_n800), .B2(new_n1120), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n287), .B2(new_n953), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G125), .C2(new_n792), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n279), .B(new_n254), .C1(new_n789), .C2(new_n1122), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G124), .B2(new_n780), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1196), .B2(new_n1200), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT117), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n835), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1190), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1171), .B2(new_n769), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1189), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1188), .A2(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1006), .B(KEYINPUT119), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1143), .A2(new_n1150), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n903), .A2(new_n768), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n759), .B1(G68), .B2(new_n836), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n790), .A2(G77), .B1(new_n805), .B2(G107), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n784), .A2(G116), .B1(new_n794), .B2(G283), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n356), .B1(new_n779), .B2(new_n842), .C1(new_n776), .C2(new_n202), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n792), .B2(G294), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1228), .A4(new_n1039), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1193), .B1(new_n1113), .B2(new_n779), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n764), .B(new_n1230), .C1(G159), .C2(new_n800), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n1068), .B2(new_n953), .C1(new_n287), .C2(new_n786), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT120), .Z(new_n1233));
  AOI22_X1  g1033(.A1(G132), .A2(new_n792), .B1(new_n784), .B2(new_n1120), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n849), .B2(new_n793), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1224), .B1(new_n1236), .B2(new_n771), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1148), .A2(new_n758), .B1(new_n1223), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1222), .A2(new_n1238), .ZN(G381));
  OR2_X1    g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  OR3_X1    g1040(.A1(G390), .A2(G384), .A3(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1241), .A2(G387), .A3(G381), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1188), .A2(new_n1217), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1105), .A2(new_n1130), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1154), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n1151), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .ZN(G407));
  INV_X1    g1047(.A(new_n1246), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n669), .A2(G213), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(G375), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT121), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1052(.A(G378), .B(new_n1217), .C1(new_n1183), .C2(new_n1187), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1186), .A2(new_n1156), .A3(new_n1221), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1189), .A2(new_n1216), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1246), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1258), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1259), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT123), .A3(new_n1219), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n687), .B1(new_n1262), .B2(KEYINPUT60), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1238), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(G384), .A3(new_n1238), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1257), .A2(new_n1249), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n669), .A2(KEYINPUT125), .A3(G213), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1270), .A2(new_n1271), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1278), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1270), .A2(new_n1271), .A3(new_n1280), .A4(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1257), .A2(new_n1249), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1257), .A2(new_n1286), .A3(new_n1249), .A4(new_n1273), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1275), .A2(new_n1284), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G393), .A2(G396), .ZN(new_n1290));
  AND3_X1   g1090(.A1(G387), .A2(new_n1240), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(G387), .A2(new_n1292), .B1(new_n1240), .B2(new_n1290), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1240), .A2(new_n1290), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G387), .ZN(new_n1296));
  AND2_X1   g1096(.A1(G387), .A2(new_n1292), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G390), .B(new_n1296), .C1(new_n1297), .C2(new_n1295), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1288), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1249), .A4(new_n1273), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1282), .A2(new_n1283), .A3(KEYINPUT126), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT126), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1274), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT124), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1274), .A2(new_n1310), .A3(new_n1307), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1300), .B1(new_n1306), .B2(new_n1312), .ZN(G405));
  OAI21_X1  g1113(.A(new_n1253), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1273), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1253), .B(new_n1272), .C1(new_n1243), .C2(new_n1248), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1315), .A2(new_n1299), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1299), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


