//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n202), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT78), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n216), .A3(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n213), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT77), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n213), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n214), .A2(KEYINPUT76), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n228), .A3(KEYINPUT2), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n219), .A2(new_n220), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n225), .A2(new_n232), .A3(new_n202), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT29), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n209), .B(KEYINPUT73), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G228gat), .A3(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G228gat), .A2(G233gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n234), .B(new_n240), .C1(new_n209), .C2(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G78gat), .B(G106gat), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT31), .B(G50gat), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT83), .ZN(new_n248));
  INV_X1    g047(.A(new_n243), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n239), .A2(new_n249), .A3(new_n241), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n248), .B1(new_n244), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(G120gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G134gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n260), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n261), .A2(new_n262), .ZN(new_n272));
  NAND2_X1  g071(.A1(G127gat), .A2(G134gat), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n258), .B2(G120gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n256), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n278), .B2(new_n257), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT71), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n233), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n254), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n224), .A2(new_n221), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n286), .A2(new_n218), .B1(new_n230), .B2(new_n231), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(new_n284), .A3(new_n271), .A4(new_n279), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n271), .A2(KEYINPUT71), .A3(new_n279), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n280), .ZN(new_n290));
  OAI211_X1 g089(.A(KEYINPUT79), .B(KEYINPUT4), .C1(new_n290), .C2(new_n233), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n202), .B1(new_n225), .B2(new_n232), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n235), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n279), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n233), .B(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n294), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(KEYINPUT5), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n284), .B(new_n287), .C1(new_n289), .C2(new_n280), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT4), .B1(new_n233), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(KEYINPUT80), .A3(new_n304), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT5), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT81), .B1(new_n309), .B2(new_n298), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n303), .A2(KEYINPUT80), .A3(new_n304), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT80), .B1(new_n303), .B2(new_n304), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n311), .B(new_n298), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n302), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT0), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G57gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G85gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT39), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n300), .A2(new_n294), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n297), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n312), .B2(new_n313), .ZN(new_n326));
  AOI211_X1 g125(.A(new_n323), .B(new_n324), .C1(new_n326), .C2(new_n294), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n323), .A3(new_n294), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT40), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(KEYINPUT84), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n327), .A2(new_n331), .B1(KEYINPUT84), .B2(new_n329), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n324), .B1(new_n326), .B2(new_n294), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT39), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n329), .A2(KEYINPUT84), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n328), .A4(new_n330), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n322), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(G64gat), .ZN(new_n339));
  INV_X1    g138(.A(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n237), .ZN(new_n343));
  INV_X1    g142(.A(G226gat), .ZN(new_n344));
  INV_X1    g143(.A(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G183gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT27), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT27), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT27), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n352), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n354), .A2(new_n359), .A3(KEYINPUT67), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT26), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n366), .B2(KEYINPUT23), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(KEYINPUT23), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n352), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT24), .A3(new_n364), .ZN(new_n379));
  AND4_X1   g178(.A1(new_n369), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT65), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n381), .A3(new_n369), .A4(new_n377), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n364), .A2(KEYINPUT24), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n380), .A2(KEYINPUT25), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(KEYINPUT25), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n373), .A2(new_n375), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(new_n377), .A3(new_n383), .A4(new_n379), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n365), .A2(new_n371), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n347), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n388), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n362), .A2(new_n371), .A3(new_n363), .A4(new_n364), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n347), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n343), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n380), .A2(new_n383), .B1(KEYINPUT25), .B2(new_n382), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n385), .A2(new_n387), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n346), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n400), .A2(new_n209), .A3(new_n393), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n342), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n395), .B2(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n210), .A3(new_n394), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n237), .B1(new_n400), .B2(new_n393), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT74), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n341), .B(KEYINPUT75), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n253), .B1(new_n337), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  INV_X1    g214(.A(new_n321), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n302), .B(new_n416), .C1(new_n310), .C2(new_n316), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n314), .B(new_n315), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n420), .B2(new_n302), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(KEYINPUT6), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n322), .A2(KEYINPUT85), .A3(new_n418), .A4(new_n417), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n409), .A3(KEYINPUT37), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n395), .B2(new_n401), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n341), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT38), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n390), .A2(new_n394), .A3(new_n343), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n209), .B1(new_n400), .B2(new_n393), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT37), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n428), .A2(new_n431), .A3(new_n410), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n402), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n414), .B1(new_n425), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n402), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(KEYINPUT38), .B2(new_n429), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(new_n423), .A3(new_n422), .A4(new_n424), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT86), .A3(new_n414), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n419), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n417), .A2(KEYINPUT82), .A3(new_n418), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n322), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n413), .B1(new_n448), .B2(new_n423), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  INV_X1    g250(.A(new_n290), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n398), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n391), .A2(new_n290), .A3(new_n392), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(G227gat), .A3(new_n454), .A4(G233gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n456));
  XNOR2_X1  g255(.A(G15gat), .B(G43gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(G71gat), .ZN(new_n458));
  INV_X1    g257(.A(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n455), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n455), .B2(new_n462), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n456), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(KEYINPUT33), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n455), .A2(KEYINPUT32), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n465), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n454), .ZN(new_n471));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n465), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT34), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n451), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n475), .A3(new_n478), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT36), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n450), .A2(new_n253), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n444), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n253), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n450), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  INV_X1    g289(.A(new_n413), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n425), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT92), .B(G57gat), .Z(new_n495));
  MUX2_X1   g294(.A(G57gat), .B(new_n495), .S(G64gat), .Z(new_n496));
  NOR2_X1   g295(.A1(G71gat), .A2(G78gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT9), .ZN(new_n498));
  NAND2_X1  g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n497), .ZN(new_n502));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n499), .B(new_n502), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT95), .B(G92gat), .ZN(new_n507));
  INV_X1    g306(.A(G85gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT8), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G99gat), .B(G106gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT96), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n513), .B(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n513), .A2(KEYINPUT99), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(KEYINPUT99), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT100), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522));
  INV_X1    g321(.A(new_n515), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n513), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n517), .B1(new_n525), .B2(new_n506), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n506), .A2(new_n516), .A3(KEYINPUT10), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT101), .ZN(new_n532));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n526), .A2(new_n533), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n529), .B1(new_n526), .B2(new_n527), .ZN(new_n536));
  INV_X1    g335(.A(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT101), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540));
  INV_X1    g339(.A(G176gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G204gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT102), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n536), .A2(new_n537), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n535), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G197gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT11), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(G169gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  INV_X1    g358(.A(G36gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT87), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR3_X1   g363(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT88), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G43gat), .B(G50gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n563), .A2(new_n565), .B1(new_n559), .B2(new_n560), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(KEYINPUT15), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n567), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT17), .ZN(new_n573));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT16), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G1gat), .ZN(new_n576));
  INV_X1    g375(.A(G8gat), .ZN(new_n577));
  OAI221_X1 g376(.A(new_n576), .B1(KEYINPUT89), .B2(new_n577), .C1(G1gat), .C2(new_n574), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT90), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n572), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT91), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n588), .A3(new_n580), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n582), .A2(new_n584), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT18), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n580), .B(new_n572), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n586), .B(KEYINPUT13), .Z(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n558), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT18), .A3(new_n587), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT18), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  AND4_X1   g398(.A1(new_n558), .A2(new_n597), .A3(new_n594), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n580), .ZN(new_n605));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n610), .A2(new_n611), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n610), .A2(new_n611), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n516), .B(KEYINPUT97), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n573), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n572), .A2(new_n516), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n262), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n629), .B(G134gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G162gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n603), .B1(new_n624), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(KEYINPUT98), .A3(new_n623), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n494), .A2(new_n553), .A3(new_n602), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n601), .B1(new_n485), .B2(new_n493), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(KEYINPUT103), .A3(new_n553), .A4(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n448), .A2(new_n423), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n413), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n575), .A2(new_n577), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n658), .A2(new_n659), .B1(G8gat), .B2(new_n657), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n663), .B2(new_n661), .ZN(G1325gat));
  NOR2_X1   g463(.A1(new_n474), .A2(new_n479), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n652), .B2(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT36), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT36), .B1(new_n481), .B2(new_n482), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n649), .B2(new_n651), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(G15gat), .B2(new_n671), .ZN(G1326gat));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n253), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT104), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n676), .A3(new_n253), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(new_n652), .B2(new_n253), .ZN(new_n679));
  AOI211_X1 g478(.A(KEYINPUT104), .B(new_n486), .C1(new_n649), .C2(new_n651), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT43), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n246), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n673), .A3(new_n677), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n679), .B2(new_n680), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(G22gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(G1327gat));
  OAI22_X1  g485(.A1(new_n667), .A2(new_n668), .B1(new_n449), .B2(new_n486), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n439), .B2(new_n443), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n490), .B1(new_n489), .B2(new_n449), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n481), .A2(new_n482), .A3(new_n490), .A4(new_n486), .ZN(new_n690));
  INV_X1    g489(.A(new_n425), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n690), .A2(new_n691), .A3(new_n413), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n642), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n640), .A2(KEYINPUT107), .A3(new_n641), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n640), .B2(new_n641), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n442), .A2(KEYINPUT86), .A3(new_n414), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT86), .B1(new_n442), .B2(new_n414), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n704), .B2(new_n687), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n444), .A2(new_n484), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n693), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n695), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n553), .A2(new_n624), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n602), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n559), .B1(new_n713), .B2(new_n654), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(new_n715), .A3(new_n642), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT105), .B1(new_n710), .B2(new_n644), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n650), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(G29gat), .A3(new_n653), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n714), .A2(new_n720), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n718), .A2(G36gat), .A3(new_n491), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n712), .B2(new_n491), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(G43gat), .B1(new_n712), .B2(new_n670), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT47), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n665), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n718), .A2(G43gat), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n726), .B(new_n730), .C1(new_n727), .C2(KEYINPUT47), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  NAND3_X1  g533(.A1(new_n713), .A2(G50gat), .A3(new_n253), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n253), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(G50gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n735), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1331gat));
  AND3_X1   g544(.A1(new_n444), .A2(new_n484), .A3(new_n706), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n706), .B1(new_n444), .B2(new_n484), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n493), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n646), .A2(new_n601), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n552), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n748), .A2(new_n752), .A3(new_n552), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n653), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n495), .ZN(G1332gat));
  NAND3_X1  g555(.A1(new_n751), .A2(new_n413), .A3(new_n753), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT49), .B(G64gat), .Z(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n754), .B2(new_n729), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n669), .A2(G71gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT50), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n762), .B(new_n766), .C1(new_n754), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n754), .A2(new_n486), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(G78gat), .Z(G1335gat));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n748), .A2(new_n700), .B1(KEYINPUT44), .B2(new_n694), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n602), .A2(new_n623), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n553), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n771), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n709), .A2(KEYINPUT111), .A3(new_n775), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n508), .B(new_n653), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n705), .A2(new_n707), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n774), .B1(new_n780), .B2(new_n493), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n781), .B2(new_n642), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n708), .A2(new_n783), .A3(new_n644), .A4(new_n774), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n654), .B(new_n552), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n779), .B1(new_n508), .B2(new_n785), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n552), .A2(new_n340), .A3(new_n413), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT112), .Z(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n782), .B2(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT113), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n788), .C1(new_n782), .C2(new_n784), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n507), .B1(new_n794), .B2(new_n413), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n784), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n709), .A2(new_n775), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n491), .ZN(new_n800));
  OAI221_X1 g599(.A(new_n797), .B1(new_n798), .B2(new_n787), .C1(new_n800), .C2(new_n507), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1337gat));
  AOI211_X1 g601(.A(new_n459), .B(new_n670), .C1(new_n777), .C2(new_n778), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n552), .B(new_n665), .C1(new_n782), .C2(new_n784), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n459), .B2(new_n804), .ZN(G1338gat));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n794), .B2(new_n253), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n806), .B(new_n552), .C1(new_n782), .C2(new_n784), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n486), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(G106gat), .B1(new_n799), .B2(new_n486), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(new_n812), .C1(new_n808), .C2(new_n486), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(new_n551), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n531), .B2(new_n533), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n548), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n534), .A2(new_n538), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .A3(new_n544), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT54), .B1(new_n534), .B2(new_n538), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n550), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n817), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n815), .B1(new_n825), .B2(KEYINPUT55), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT114), .B1(new_n820), .B2(new_n544), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n823), .A2(new_n822), .A3(new_n550), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n827), .A2(new_n828), .B1(new_n548), .B2(new_n816), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n831), .A3(new_n602), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n591), .A2(new_n558), .A3(new_n594), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n592), .A2(new_n593), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n596), .B2(new_n587), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n557), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n547), .B2(new_n551), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n698), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n837), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n698), .A2(new_n826), .A3(new_n831), .A4(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n624), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g643(.A1(new_n553), .A2(new_n643), .A3(new_n645), .A4(new_n601), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n487), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n653), .A2(new_n413), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n601), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n258), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n553), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n256), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n849), .A2(new_n624), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n268), .A2(new_n269), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n263), .A2(new_n265), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n847), .A2(new_n857), .A3(new_n642), .A4(new_n848), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n849), .B2(new_n644), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n864), .A3(new_n860), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n846), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n253), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n601), .B1(new_n829), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n838), .B1(new_n871), .B2(new_n826), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n842), .B1(new_n872), .B2(new_n642), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n845), .B1(new_n873), .B2(new_n624), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT57), .B1(new_n874), .B2(new_n486), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n670), .A2(new_n848), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT116), .Z(new_n877));
  INV_X1    g676(.A(G141gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n601), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n869), .A2(new_n875), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n876), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n867), .A2(new_n253), .A3(new_n602), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n878), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT58), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n880), .A2(new_n883), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n880), .C2(new_n883), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n885), .A2(new_n886), .B1(new_n890), .B2(new_n891), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n867), .A2(new_n253), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n876), .ZN(new_n894));
  INV_X1    g693(.A(G148gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n552), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n486), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n845), .B(KEYINPUT120), .Z(new_n900));
  NAND4_X1  g699(.A1(new_n826), .A2(new_n831), .A3(new_n642), .A4(new_n841), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n872), .B2(new_n642), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n904), .B(new_n901), .C1(new_n872), .C2(new_n642), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n624), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n868), .B1(new_n867), .B2(new_n253), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n908), .A2(new_n552), .A3(new_n877), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n897), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n869), .A2(new_n875), .A3(new_n877), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n897), .B1(new_n913), .B2(new_n553), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n895), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n896), .B1(new_n912), .B2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n913), .B2(new_n624), .ZN(new_n917));
  INV_X1    g716(.A(G155gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n918), .A3(new_n623), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1346gat));
  NAND4_X1  g719(.A1(new_n869), .A2(new_n875), .A3(new_n698), .A4(new_n877), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n644), .A2(G162gat), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n921), .A2(G162gat), .B1(new_n894), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n654), .A2(new_n491), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n847), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n601), .ZN(new_n927));
  XNOR2_X1  g726(.A(KEYINPUT123), .B(G169gat), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(G1348gat));
  NOR2_X1   g728(.A1(new_n926), .A2(new_n553), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(new_n541), .ZN(G1349gat));
  OAI21_X1  g730(.A(new_n348), .B1(new_n926), .B2(new_n624), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n349), .A2(new_n351), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n847), .A2(new_n933), .A3(new_n623), .A4(new_n925), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g735(.A1(new_n847), .A2(new_n642), .A3(new_n925), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n847), .A2(new_n352), .A3(new_n698), .A4(new_n925), .ZN(new_n946));
  NAND2_X1  g745(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n940), .A2(new_n941), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(G1351gat));
  NAND2_X1  g749(.A1(new_n670), .A2(new_n925), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n907), .A2(new_n909), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n602), .ZN(new_n953));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n654), .B1(new_n844), .B2(new_n846), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n670), .A2(new_n413), .A3(new_n253), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n602), .A2(new_n954), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n953), .A2(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NOR3_X1   g759(.A1(new_n958), .A2(G204gat), .A3(new_n553), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT62), .ZN(new_n962));
  NOR4_X1   g761(.A1(new_n907), .A2(new_n909), .A3(new_n553), .A4(new_n951), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n543), .B2(new_n963), .ZN(G1353gat));
  NOR4_X1   g763(.A1(new_n907), .A2(new_n909), .A3(new_n624), .A4(new_n951), .ZN(new_n965));
  OAI211_X1 g764(.A(KEYINPUT127), .B(KEYINPUT63), .C1(new_n965), .C2(new_n204), .ZN(new_n966));
  INV_X1    g765(.A(new_n951), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n908), .A2(new_n623), .A3(new_n910), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g767(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n969));
  NAND2_X1  g768(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n968), .A2(G211gat), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n204), .A3(new_n623), .A4(new_n957), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(G1354gat));
  NOR2_X1   g772(.A1(new_n644), .A2(new_n205), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n955), .A2(new_n698), .A3(new_n957), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n952), .A2(new_n974), .B1(new_n205), .B2(new_n975), .ZN(G1355gat));
endmodule


