//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n208), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n208), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n216), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n203), .A2(new_n205), .ZN(new_n230));
  INV_X1    g0030(.A(G50), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n232), .A2(G20), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n236));
  NAND4_X1  g0036(.A1(new_n218), .A2(new_n229), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n201), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT66), .B(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND2_X1  g0055(.A1(new_n209), .A2(G45), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT5), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT5), .A2(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT81), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G274), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  INV_X1    g0063(.A(new_n258), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT5), .A2(G41), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n263), .B(G274), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT81), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n261), .A2(new_n267), .B1(new_n271), .B2(G270), .ZN(new_n272));
  INV_X1    g0072(.A(G303), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT68), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n273), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT75), .B1(new_n274), .B2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT75), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n276), .A3(KEYINPUT3), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(new_n280), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n216), .A2(G1698), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G257), .B2(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n270), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n272), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT85), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n272), .A2(new_n291), .A3(KEYINPUT85), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G116), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n233), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n276), .A2(G1), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n297), .B1(new_n303), .B2(G116), .ZN(new_n304));
  AOI21_X1  g0104(.A(G20), .B1(G33), .B2(G283), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n276), .A2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT86), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT86), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G116), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n298), .A2(new_n233), .B1(G20), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(KEYINPUT20), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT20), .B1(new_n311), .B2(new_n313), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n304), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n294), .A2(new_n295), .A3(G169), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT21), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n272), .A2(new_n291), .A3(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n317), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  INV_X1    g0123(.A(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n325), .B2(new_n304), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n326), .A2(KEYINPUT21), .A3(new_n294), .A4(new_n295), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n295), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT85), .B1(new_n272), .B2(new_n291), .ZN(new_n330));
  OAI21_X1  g0130(.A(G190), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n317), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n294), .A2(G200), .A3(new_n295), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n210), .B1(new_n230), .B2(new_n231), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n210), .A2(G33), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G20), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n299), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n209), .A2(G20), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G50), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n343), .B1(G50), .B2(new_n296), .C1(new_n301), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n209), .A2(G274), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT67), .B(G45), .Z(new_n348));
  INV_X1    g0148(.A(G41), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n269), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n281), .B1(new_n279), .B2(new_n280), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G1698), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G222), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(G223), .A3(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n224), .C2(new_n358), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n355), .B1(new_n362), .B2(new_n270), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n346), .B1(new_n363), .B2(G169), .ZN(new_n364));
  INV_X1    g0164(.A(G179), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n346), .B1(KEYINPUT69), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n363), .A2(G190), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n370), .A2(new_n376), .A3(new_n372), .A4(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n366), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n296), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n299), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(G77), .A3(new_n344), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G77), .B2(new_n296), .ZN(new_n382));
  INV_X1    g0182(.A(new_n337), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n340), .B1(G20), .B2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n338), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n299), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n270), .B1(new_n358), .B2(G107), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n278), .A2(new_n282), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G232), .A2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n220), .B2(G1698), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n351), .B1(new_n225), .B2(new_n354), .C1(new_n388), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(new_n393), .B2(new_n323), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n387), .C1(new_n397), .C2(new_n393), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n378), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  INV_X1    g0201(.A(G232), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n354), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n269), .A2(new_n353), .A3(KEYINPUT78), .A4(G232), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n350), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n352), .A2(G1698), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G223), .B2(G1698), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n287), .A2(new_n407), .B1(new_n276), .B2(new_n221), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n270), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(G190), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n415), .B2(new_n371), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n383), .A2(new_n344), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n417), .A2(new_n301), .B1(new_n296), .B2(new_n383), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT3), .B(G33), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(G20), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n420), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(KEYINPUT76), .B(new_n423), .C1(new_n275), .C2(new_n277), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(G20), .B1(new_n278), .B2(new_n282), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G68), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(G20), .B1(G159), .B2(new_n340), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n287), .A2(new_n422), .A3(new_n210), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n422), .B1(new_n287), .B2(new_n210), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT16), .B(new_n432), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n299), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n419), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n400), .B1(new_n416), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT16), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n210), .B1(new_n356), .B2(new_n357), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n202), .ZN(new_n444));
  INV_X1    g0244(.A(new_n432), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n438), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n418), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n409), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT79), .B1(new_n405), .B2(new_n409), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n371), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n411), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n440), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n439), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n410), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n415), .A2(new_n323), .B1(new_n365), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT77), .B(new_n419), .C1(new_n433), .C2(new_n438), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n455), .B1(KEYINPUT18), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n457), .A2(new_n463), .A3(new_n459), .A4(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT80), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n379), .A2(new_n202), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT12), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n380), .A2(G68), .A3(new_n344), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT11), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n341), .A2(new_n231), .B1(new_n210), .B2(G68), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n338), .A2(new_n224), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n299), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n469), .B2(new_n472), .ZN(new_n474));
  XOR2_X1   g0274(.A(new_n474), .B(KEYINPUT72), .Z(new_n475));
  INV_X1    g0275(.A(KEYINPUT14), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT13), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n402), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G226), .B2(G1698), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n356), .A2(new_n357), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n270), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT67), .B(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G41), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n485), .A2(new_n347), .B1(new_n220), .B2(new_n354), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n477), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G226), .A2(G1698), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n402), .B2(G1698), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n278), .A2(new_n282), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n269), .B1(new_n491), .B2(new_n481), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(KEYINPUT13), .A3(new_n486), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n476), .B(G169), .C1(new_n488), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n481), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n486), .B1(new_n497), .B2(new_n270), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n477), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT13), .B1(new_n492), .B2(new_n486), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT73), .A3(new_n476), .A4(G169), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT74), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT70), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n498), .B2(new_n477), .ZN(new_n506));
  NOR4_X1   g0306(.A1(new_n492), .A2(new_n486), .A3(KEYINPUT70), .A4(KEYINPUT13), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n488), .A2(new_n365), .ZN(new_n509));
  OAI21_X1  g0309(.A(G169), .B1(new_n488), .B2(new_n493), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(KEYINPUT14), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n503), .A2(new_n504), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n504), .B1(new_n503), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n475), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n488), .A2(new_n397), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT71), .ZN(new_n517));
  INV_X1    g0317(.A(new_n475), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n501), .A2(G200), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n399), .A2(new_n465), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n462), .A2(KEYINPUT80), .A3(new_n464), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n215), .A2(G1698), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G250), .B2(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n287), .A2(new_n528), .B1(new_n276), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n270), .B1(new_n271), .B2(G264), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n261), .A2(new_n267), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n323), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n270), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n271), .A2(G264), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n526), .A2(new_n533), .B1(new_n537), .B2(G179), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT87), .B1(new_n537), .B2(new_n323), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n221), .A2(KEYINPUT22), .A3(G20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n358), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n284), .A2(new_n286), .A3(new_n210), .A4(new_n280), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT22), .B1(new_n543), .B2(new_n221), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT23), .B1(new_n226), .B2(G20), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n540), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n551), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT24), .B(new_n553), .C1(new_n542), .C2(new_n544), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n299), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT25), .B1(new_n379), .B2(new_n226), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n379), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n303), .A2(G107), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n538), .A2(new_n539), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n536), .A2(new_n371), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G190), .B2(new_n536), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n269), .A2(G250), .A3(new_n256), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n209), .A2(G45), .A3(G274), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT82), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n225), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G238), .B2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n546), .B1(new_n287), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n270), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  INV_X1    g0378(.A(new_n385), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n296), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  INV_X1    g0381(.A(G97), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n338), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n482), .A2(KEYINPUT19), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT83), .B1(new_n584), .B2(new_n210), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT83), .B(new_n210), .C1(new_n481), .C2(new_n581), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n221), .A2(new_n582), .A3(new_n226), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI221_X1 g0388(.A(new_n583), .B1(new_n543), .B2(new_n202), .C1(new_n585), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n580), .B1(new_n589), .B2(new_n299), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n380), .B1(G1), .B2(new_n276), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n221), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n303), .A2(KEYINPUT84), .A3(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n572), .A2(G190), .A3(new_n576), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n578), .A2(new_n590), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n577), .A2(new_n323), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n585), .A2(new_n588), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n583), .B1(new_n543), .B2(new_n202), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n299), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n580), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n303), .A2(new_n579), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n572), .A2(new_n365), .A3(new_n576), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT4), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n225), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n278), .A2(new_n359), .A3(new_n282), .A4(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n278), .A2(G250), .A3(G1698), .A4(new_n282), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n359), .A2(G244), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n287), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G33), .A2(G283), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n610), .A2(new_n611), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n270), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n271), .A2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n532), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n270), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G190), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n443), .A2(new_n226), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT6), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n625), .A2(new_n582), .A3(G107), .ZN(new_n626));
  XNOR2_X1  g0426(.A(G97), .B(G107), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n628), .A2(new_n210), .B1(new_n224), .B2(new_n341), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n299), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n296), .A2(G97), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n303), .B2(G97), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n621), .A2(new_n623), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n620), .A2(new_n323), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n629), .B1(new_n429), .B2(G107), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n300), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n622), .A2(new_n365), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n607), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n335), .A2(new_n525), .A3(new_n565), .A4(new_n639), .ZN(G372));
  AND2_X1   g0440(.A1(new_n440), .A2(new_n454), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT88), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n395), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n394), .B(KEYINPUT88), .C1(G179), .C2(new_n393), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n520), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n514), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n459), .A2(new_n439), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(new_n463), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n375), .A2(new_n377), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n366), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n639), .B(new_n563), .C1(new_n328), .C2(new_n560), .ZN(new_n654));
  INV_X1    g0454(.A(new_n606), .ZN(new_n655));
  INV_X1    g0455(.A(new_n638), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n607), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n597), .A2(new_n606), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n638), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n653), .B1(new_n524), .B2(new_n662), .ZN(G369));
  NAND3_X1  g0463(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n335), .B1(new_n332), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n328), .A2(new_n317), .A3(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(KEYINPUT90), .A3(new_n676), .ZN(new_n680));
  INV_X1    g0480(.A(new_n560), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n563), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n670), .B1(new_n555), .B2(new_n559), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n681), .B2(new_n670), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n679), .A2(new_n680), .A3(G330), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n328), .A2(new_n670), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n681), .A2(new_n669), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(G399));
  OAI21_X1  g0490(.A(KEYINPUT91), .B1(new_n214), .B2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n214), .A2(KEYINPUT91), .A3(G41), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n587), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n232), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n697), .B(KEYINPUT92), .C1(new_n698), .C2(new_n695), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(KEYINPUT92), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT28), .Z(new_n701));
  AOI21_X1  g0501(.A(new_n669), .B1(new_n654), .B2(new_n661), .ZN(new_n702));
  AND2_X1   g0502(.A1(KEYINPUT93), .A2(KEYINPUT29), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(KEYINPUT93), .A2(KEYINPUT29), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n702), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n531), .A2(new_n576), .A3(new_n572), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n321), .A2(new_n709), .A3(new_n622), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n577), .A2(new_n365), .A3(new_n536), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n294), .A3(new_n295), .A4(new_n620), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n321), .A2(new_n709), .A3(new_n622), .A4(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n669), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n335), .A2(new_n565), .A3(new_n639), .A4(new_n670), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n708), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n707), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n701), .B1(new_n727), .B2(G1), .ZN(G364));
  NAND2_X1  g0528(.A1(new_n679), .A2(new_n680), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n708), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n679), .A2(new_n680), .A3(G330), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n210), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n209), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n694), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  INV_X1    g0538(.A(new_n287), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n214), .A2(new_n739), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n740), .B1(new_n698), .B2(new_n484), .C1(new_n251), .C2(new_n262), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n358), .A2(new_n213), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n743), .A2(G355), .B1(new_n312), .B2(new_n214), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n233), .B1(G20), .B2(new_n323), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(new_n365), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n753), .A2(new_n371), .A3(G190), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n753), .A2(new_n397), .A3(G200), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(G322), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n397), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n397), .A2(new_n371), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n758), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G283), .A2(new_n760), .B1(new_n763), .B2(G303), .ZN(new_n764));
  INV_X1    g0564(.A(G329), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n757), .B(new_n764), .C1(new_n765), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n761), .A2(new_n752), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n752), .A2(new_n766), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G326), .A2(new_n773), .B1(new_n775), .B2(G311), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n397), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n210), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n389), .C1(new_n529), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n754), .A2(G68), .B1(new_n773), .B2(G50), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n760), .A2(G107), .B1(new_n775), .B2(G77), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n756), .A2(G58), .B1(G87), .B2(new_n763), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n358), .C1(new_n582), .C2(new_n778), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n771), .A2(new_n779), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n736), .B1(new_n788), .B2(new_n749), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n751), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n677), .B2(new_n748), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n738), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n387), .A2(new_n670), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n643), .A2(new_n644), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n395), .B(new_n398), .C1(new_n387), .C2(new_n670), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n702), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n724), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n735), .B1(new_n799), .B2(new_n724), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(KEYINPUT98), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT98), .B2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(new_n749), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n747), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n735), .B1(G77), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n756), .A2(G143), .B1(new_n773), .B2(G137), .ZN(new_n807));
  INV_X1    g0607(.A(new_n754), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n339), .B2(new_n808), .C1(new_n780), .C2(new_n774), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  INV_X1    g0610(.A(new_n770), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G132), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n759), .A2(new_n202), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n287), .B(new_n813), .C1(G50), .C2(new_n763), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(new_n201), .C2(new_n778), .ZN(new_n815));
  INV_X1    g0615(.A(new_n756), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(new_n529), .B1(new_n582), .B2(new_n778), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n759), .A2(new_n221), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n772), .A2(new_n273), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G283), .C2(new_n754), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n811), .A2(G311), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G116), .A2(new_n775), .B1(new_n763), .B2(G107), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n821), .A2(new_n822), .A3(new_n389), .A4(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n810), .A2(new_n815), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n806), .B1(new_n825), .B2(new_n749), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n797), .B2(new_n747), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n803), .A2(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT35), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n628), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n830), .A2(G20), .A3(G116), .A4(new_n234), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT99), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(new_n829), .B2(new_n628), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n835));
  XNOR2_X1  g0635(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n232), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n231), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n209), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT37), .B1(new_n448), .B2(new_n453), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n461), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT101), .ZN(new_n844));
  INV_X1    g0644(.A(new_n667), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n457), .A2(new_n844), .A3(new_n460), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n457), .A2(new_n460), .A3(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n843), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n846), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT102), .B1(new_n416), .B2(new_n439), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n448), .A2(new_n453), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n853), .A3(new_n649), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT103), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n851), .A2(new_n853), .A3(new_n856), .A4(new_n649), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n850), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n849), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n850), .B1(new_n641), .B2(new_n650), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n841), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n461), .A2(KEYINPUT18), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n641), .A2(new_n862), .A3(new_n464), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n441), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n419), .B1(new_n865), .B2(new_n438), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n845), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n459), .A2(new_n866), .B1(new_n448), .B2(new_n453), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n867), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(KEYINPUT38), .C1(new_n872), .C2(new_n849), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT39), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n867), .B1(new_n462), .B2(new_n464), .ZN(new_n875));
  INV_X1    g0675(.A(new_n843), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n850), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n841), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n514), .A2(new_n669), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n702), .A2(new_n797), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n395), .B2(new_n669), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n475), .A2(new_n669), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n514), .A2(new_n520), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n475), .B(new_n669), .C1(new_n512), .C2(new_n513), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n873), .B2(new_n878), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n650), .A2(new_n845), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n522), .A2(new_n706), .A3(new_n523), .A4(new_n704), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n653), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n524), .B1(new_n723), .B2(new_n722), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n798), .B1(new_n722), .B2(new_n723), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n861), .B2(new_n873), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n878), .A2(new_n873), .ZN(new_n901));
  AND4_X1   g0701(.A1(new_n335), .A2(new_n639), .A3(new_n565), .A4(new_n670), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n797), .B1(new_n902), .B2(new_n721), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n886), .B2(new_n887), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n708), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n897), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n209), .B2(new_n732), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n896), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n840), .B1(new_n910), .B2(new_n911), .ZN(G367));
  NAND2_X1  g0712(.A1(new_n636), .A2(new_n669), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n633), .A2(new_n638), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n638), .B2(new_n670), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n638), .B1(new_n919), .B2(new_n681), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n670), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n917), .A2(new_n918), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n687), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT105), .ZN(new_n924));
  INV_X1    g0724(.A(new_n687), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n923), .A2(KEYINPUT42), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT42), .B1(new_n923), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n670), .B1(new_n590), .B2(new_n595), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n655), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n659), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT106), .B1(new_n929), .B2(new_n934), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n685), .A2(new_n919), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n935), .A2(new_n938), .A3(new_n940), .A4(new_n937), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n694), .B(KEYINPUT41), .Z(new_n944));
  INV_X1    g0744(.A(new_n686), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n684), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n731), .A2(new_n925), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n925), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n679), .A2(new_n680), .A3(G330), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n726), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT44), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n922), .B2(new_n689), .ZN(new_n952));
  INV_X1    g0752(.A(new_n689), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(KEYINPUT44), .A3(new_n919), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n922), .A2(KEYINPUT45), .A3(new_n689), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n953), .B2(new_n919), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n685), .B1(new_n961), .B2(KEYINPUT107), .ZN(new_n962));
  INV_X1    g0762(.A(new_n685), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n960), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n950), .B(new_n962), .C1(KEYINPUT107), .C2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n944), .B1(new_n965), .B2(new_n727), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n942), .B(new_n943), .C1(new_n966), .C2(new_n734), .ZN(new_n967));
  INV_X1    g0767(.A(new_n740), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n750), .B1(new_n213), .B2(new_n385), .C1(new_n968), .C2(new_n246), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n735), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n748), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n816), .A2(new_n273), .ZN(new_n972));
  INV_X1    g0772(.A(new_n767), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n739), .B(new_n972), .C1(G317), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n778), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G107), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n763), .A2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n759), .A2(new_n582), .ZN(new_n979));
  INV_X1    g0779(.A(G311), .ZN(new_n980));
  INV_X1    g0780(.A(G283), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n772), .A2(new_n980), .B1(new_n774), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n979), .B(new_n982), .C1(G294), .C2(new_n754), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n974), .A2(new_n976), .A3(new_n978), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n975), .A2(G68), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n773), .A2(G143), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n816), .C2(new_n339), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT108), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n358), .B1(new_n224), .B2(new_n759), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G58), .A2(new_n763), .B1(new_n973), .B2(G137), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n754), .A2(G159), .B1(G50), .B2(new_n775), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n984), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n970), .B1(new_n971), .B2(new_n932), .C1(new_n998), .C2(new_n804), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n967), .A2(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n950), .A2(new_n695), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n947), .A2(new_n949), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n727), .B2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n684), .A2(new_n971), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n383), .A2(new_n231), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT50), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n696), .B(new_n262), .C1(new_n202), .C2(new_n224), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n740), .B1(new_n1006), .B2(new_n1007), .C1(new_n243), .C2(new_n348), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n743), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(G107), .B2(new_n213), .C1(new_n696), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT111), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n750), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n754), .A2(new_n383), .B1(G68), .B2(new_n775), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT112), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n762), .A2(new_n224), .B1(new_n767), .B2(new_n339), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G50), .B2(new_n756), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n780), .A2(new_n772), .B1(new_n759), .B2(new_n582), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n287), .B(new_n1019), .C1(new_n579), .C2(new_n975), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n760), .A2(G116), .B1(new_n973), .B2(G326), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n778), .A2(new_n981), .B1(new_n762), .B2(new_n529), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n756), .A2(G317), .B1(new_n773), .B2(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n273), .B2(new_n774), .C1(new_n980), .C2(new_n808), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n287), .B(new_n1022), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1021), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n736), .B(new_n1014), .C1(new_n749), .C2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1002), .A2(new_n734), .B1(new_n1004), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1003), .A2(new_n1034), .ZN(G393));
  XNOR2_X1  g0835(.A(new_n960), .B(new_n685), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n965), .B(new_n694), .C1(new_n950), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n919), .A2(new_n748), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n750), .B1(new_n582), .B2(new_n213), .C1(new_n968), .C2(new_n254), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n735), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n808), .A2(new_n273), .B1(new_n759), .B2(new_n226), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n358), .B(new_n1041), .C1(G116), .C2(new_n975), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n775), .B1(new_n973), .B2(G322), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n981), .C2(new_n762), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n756), .A2(G311), .B1(new_n773), .B2(G317), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n756), .A2(G159), .B1(new_n773), .B2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n287), .B(new_n819), .C1(G143), .C2(new_n973), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n754), .A2(G50), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n383), .A2(new_n775), .B1(new_n763), .B2(G68), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n975), .A2(G77), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1044), .A2(new_n1046), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1040), .B1(new_n1054), .B2(new_n749), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1036), .A2(new_n734), .B1(new_n1038), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1037), .A2(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(new_n881), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n889), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n874), .B2(new_n879), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n861), .A2(new_n873), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n1058), .A3(new_n889), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n888), .A2(new_n898), .A3(G330), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1064), .A3(new_n1062), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n734), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n522), .A2(new_n523), .A3(new_n724), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n894), .A2(new_n653), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n888), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n724), .A2(KEYINPUT113), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n797), .B1(new_n724), .B2(KEYINPUT113), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n884), .B1(new_n1077), .B2(new_n1064), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n708), .B2(new_n903), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1079), .A2(new_n1064), .A3(new_n884), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1073), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1071), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n694), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n735), .B1(new_n383), .B2(new_n805), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n816), .A2(new_n312), .B1(new_n772), .B2(new_n981), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n808), .A2(new_n226), .B1(new_n774), .B2(new_n582), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n813), .B(new_n358), .C1(G87), .C2(new_n763), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n811), .A2(G294), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1089), .A2(new_n1052), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n763), .A2(G150), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1093), .A2(KEYINPUT53), .B1(new_n780), .B2(new_n778), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n389), .B(new_n1094), .C1(KEYINPUT53), .C2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n811), .A2(G125), .ZN(new_n1096));
  INV_X1    g0896(.A(G137), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n808), .A2(new_n1097), .B1(new_n759), .B2(new_n231), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n775), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n756), .A2(G132), .B1(new_n773), .B2(G128), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT115), .Z(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT116), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n804), .B1(new_n1105), .B2(KEYINPUT116), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1086), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n880), .B2(new_n747), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1070), .A2(new_n1085), .A3(new_n1109), .ZN(G378));
  NAND2_X1  g0910(.A1(new_n346), .A2(new_n845), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n378), .B(new_n1111), .Z(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n746), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n735), .B1(G50), .B2(new_n805), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n739), .A2(G33), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G50), .B1(new_n1118), .B2(new_n349), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT117), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G116), .A2(new_n773), .B1(new_n760), .B2(G58), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n226), .B2(new_n816), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G283), .B2(new_n811), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n754), .A2(G97), .B1(new_n579), .B2(new_n775), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT118), .ZN(new_n1125));
  AOI211_X1 g0925(.A(G41), .B(new_n739), .C1(G77), .C2(new_n763), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1125), .A3(new_n985), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1120), .B1(new_n1128), .B2(KEYINPUT58), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n276), .B(new_n349), .C1(new_n759), .C2(new_n780), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G124), .B2(new_n973), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n754), .A2(G132), .B1(new_n773), .B2(G125), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n816), .C1(new_n1097), .C2(new_n774), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n763), .A2(KEYINPUT119), .A3(new_n1100), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n762), .B2(new_n1099), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n339), .C2(new_n778), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT120), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1131), .B1(new_n1141), .B2(KEYINPUT59), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT59), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1129), .B1(KEYINPUT58), .B2(new_n1128), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT121), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n804), .B1(new_n1145), .B2(KEYINPUT121), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1117), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1116), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n888), .A2(new_n898), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n873), .B2(new_n878), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n1152), .B2(KEYINPUT40), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT122), .B1(new_n1153), .B2(new_n900), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n901), .A2(new_n904), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT40), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n708), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT122), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n900), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1114), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n1115), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n893), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n900), .A2(new_n905), .A3(KEYINPUT122), .A4(new_n708), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1115), .B1(new_n1165), .B2(new_n1162), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n882), .A2(new_n892), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1154), .A2(new_n1114), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n1170), .B2(new_n734), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1073), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1164), .A2(new_n1169), .B1(new_n1172), .B2(new_n1084), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n694), .B1(new_n1173), .B2(KEYINPUT57), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT123), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1164), .A2(new_n1175), .A3(new_n1169), .ZN(new_n1176));
  OAI211_X1 g0976(.A(KEYINPUT123), .B(new_n893), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1084), .B2(new_n1172), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1171), .B1(new_n1174), .B2(new_n1180), .ZN(G375));
  INV_X1    g0981(.A(new_n944), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1073), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1082), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1078), .A2(new_n733), .A3(new_n1080), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1074), .A2(new_n746), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n735), .B1(G68), .B2(new_n805), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G77), .A2(new_n760), .B1(new_n763), .B2(G97), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n389), .C1(new_n385), .C2(new_n778), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n756), .A2(G283), .B1(G107), .B2(new_n775), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n754), .A2(G116), .B1(new_n773), .B2(G294), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n770), .C2(new_n273), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n756), .A2(G137), .B1(G150), .B2(new_n775), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n754), .A2(new_n1100), .B1(new_n773), .B2(G132), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n770), .C2(new_n1133), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G58), .A2(new_n760), .B1(new_n763), .B2(G159), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n739), .C1(new_n231), .C2(new_n778), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1189), .A2(new_n1192), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1187), .B1(new_n1198), .B2(new_n749), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1185), .B1(new_n1186), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1184), .A2(new_n1200), .ZN(G381));
  XNOR2_X1  g1001(.A(G375), .B(KEYINPUT124), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1070), .A2(new_n1085), .A3(new_n1109), .ZN(new_n1203));
  INV_X1    g1003(.A(G390), .ZN(new_n1204));
  INV_X1    g1004(.A(G384), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n792), .A2(new_n1003), .A3(new_n1034), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1206), .A2(G387), .A3(G381), .A4(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1202), .A2(new_n1203), .A3(new_n1208), .ZN(G407));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G343), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1202), .A2(new_n1203), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(G407), .A2(new_n1212), .A3(G213), .ZN(G409));
  OAI211_X1 g1013(.A(G378), .B(new_n1171), .C1(new_n1174), .C2(new_n1180), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1176), .A2(new_n734), .A3(new_n1177), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1084), .A2(new_n1172), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1161), .A2(new_n1163), .A3(new_n893), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1182), .B(new_n1217), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1149), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1203), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1214), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1211), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1183), .B1(new_n1081), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1073), .B(KEYINPUT60), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n694), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1229), .A2(G384), .A3(new_n1200), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1229), .B2(new_n1200), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1223), .A2(new_n1224), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1211), .B1(new_n1214), .B2(new_n1222), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1232), .ZN(new_n1238));
  INV_X1    g1038(.A(G2897), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1224), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1232), .A2(KEYINPUT125), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1229), .A2(new_n1200), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1205), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1229), .A2(G384), .A3(new_n1200), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT125), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1239), .B2(new_n1224), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1241), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1150), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G378), .B1(new_n1251), .B2(new_n1215), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1170), .A2(new_n734), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1149), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1170), .A2(new_n1217), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n695), .B1(new_n1255), .B2(new_n1178), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1252), .B1(new_n1258), .B2(G378), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1250), .B1(new_n1259), .B2(new_n1211), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1234), .A2(new_n1235), .A3(new_n1238), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1204), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n967), .A2(G390), .A3(new_n999), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G396), .A2(G393), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1207), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n967), .B2(new_n999), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1262), .A2(new_n1268), .A3(new_n1263), .A4(new_n1266), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1261), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1274));
  AND4_X1   g1074(.A1(KEYINPUT125), .A2(new_n1243), .A3(new_n1244), .A4(new_n1240), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1240), .B1(new_n1232), .B2(KEYINPUT125), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1248), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1274), .B(new_n1235), .C1(new_n1236), .C2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT127), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1233), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1233), .A2(new_n1281), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1236), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1232), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1273), .A2(new_n1285), .ZN(G405));
  INV_X1    g1086(.A(new_n1214), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1258), .A2(G378), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1272), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1274), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1289), .A2(new_n1291), .A3(new_n1232), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1232), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G402));
endmodule


