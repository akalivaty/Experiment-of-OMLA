//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT29), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT71), .B(KEYINPUT22), .Z(new_n212));
  OAI211_X1 g011(.A(new_n206), .B(new_n207), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n218), .B2(new_n208), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n219), .B2(new_n206), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n205), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G141gat), .B(G148gat), .Z(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT77), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G155gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT77), .B(G155gat), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT78), .B(KEYINPUT2), .C1(new_n236), .C2(new_n228), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n225), .B1(new_n224), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n244));
  INV_X1    g043(.A(new_n207), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n213), .ZN(new_n247));
  INV_X1    g046(.A(new_n240), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n235), .A2(new_n237), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n222), .B(new_n248), .C1(new_n249), .C2(new_n226), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n205), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n247), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n238), .A2(KEYINPUT3), .A3(new_n240), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(KEYINPUT29), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT84), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n204), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n204), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(new_n247), .B2(new_n205), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(new_n241), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT85), .B1(new_n261), .B2(new_n251), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n204), .B1(new_n223), .B2(new_n242), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G22gat), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n258), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n258), .B2(new_n266), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(G50gat), .Z(new_n271));
  NOR3_X1   g070(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n261), .A2(new_n251), .A3(KEYINPUT85), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n264), .B1(new_n263), .B2(new_n256), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n256), .A2(KEYINPUT84), .B1(new_n242), .B2(new_n223), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n251), .A2(new_n252), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n259), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(G22gat), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n266), .A3(new_n267), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n203), .B1(new_n272), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n271), .B1(new_n268), .B2(new_n269), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n273), .A3(new_n281), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n202), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G127gat), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G134gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT1), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT68), .B(G120gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(G113gat), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT69), .B1(new_n297), .B2(G113gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n293), .B2(G113gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n296), .A2(new_n300), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n311), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n309), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n310), .A2(KEYINPUT64), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n317), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT65), .B1(new_n325), .B2(KEYINPUT25), .ZN(new_n326));
  AND2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  OR2_X1    g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n315), .ZN(new_n329));
  INV_X1    g128(.A(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n308), .C1(new_n310), .C2(KEYINPUT64), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n320), .A2(KEYINPUT64), .A3(new_n321), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n313), .B(new_n329), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n318), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n319), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(KEYINPUT27), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G183gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n341), .A3(new_n331), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT27), .B(G183gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n312), .A2(KEYINPUT26), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n314), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n348), .B(new_n320), .C1(new_n350), .C2(new_n312), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT66), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n344), .B2(new_n346), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT66), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n307), .B1(new_n338), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n319), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n320), .A2(new_n321), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT64), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(new_n324), .A3(new_n332), .A4(new_n308), .ZN(new_n364));
  INV_X1    g163(.A(new_n317), .ZN(new_n365));
  AOI211_X1 g164(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n336), .B1(new_n335), .B2(new_n318), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n306), .A2(new_n302), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n292), .A2(new_n295), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n299), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n347), .A2(KEYINPUT66), .A3(new_n352), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT66), .B1(new_n347), .B2(new_n352), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G227gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n376), .A2(new_n380), .B1(KEYINPUT70), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n375), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT32), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G15gat), .B(G43gat), .Z(new_n388));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n381), .A2(KEYINPUT70), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n390), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n384), .B(KEYINPUT32), .C1(new_n386), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n391), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n383), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n382), .A3(new_n396), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n283), .A2(new_n286), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n371), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n369), .B(KEYINPUT79), .C1(new_n299), .C2(new_n370), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n238), .B2(new_n240), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n250), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n241), .A2(new_n307), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n241), .A2(new_n307), .A3(KEYINPUT4), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n408), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n405), .A2(new_n406), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n409), .B1(new_n418), .B2(new_n241), .ZN(new_n419));
  INV_X1    g218(.A(new_n413), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR4_X1   g220(.A1(new_n371), .A2(new_n238), .A3(new_n410), .A4(new_n240), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT4), .B1(new_n241), .B2(new_n307), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n413), .A4(new_n408), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT81), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT81), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n408), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(G57gat), .B(G85gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n426), .A2(new_n431), .A3(new_n436), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n403), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n205), .B(new_n445), .C1(new_n338), .C2(new_n356), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n368), .A2(new_n447), .A3(new_n374), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n254), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n368), .B2(new_n353), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT29), .B1(new_n368), .B2(new_n374), .ZN(new_n452));
  OAI22_X1  g251(.A1(new_n450), .A2(new_n451), .B1(new_n452), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n205), .B1(new_n338), .B2(new_n358), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n445), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n247), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n447), .B1(new_n338), .B2(new_n356), .ZN(new_n459));
  AOI22_X1  g258(.A1(KEYINPUT73), .A2(new_n459), .B1(new_n454), .B2(new_n445), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n452), .A2(new_n450), .A3(new_n447), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n254), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT74), .ZN(new_n463));
  XOR2_X1   g262(.A(G8gat), .B(G36gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT75), .ZN(new_n465));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n458), .A2(KEYINPUT30), .A3(new_n463), .A4(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n457), .B(new_n254), .C1(new_n460), .C2(new_n461), .ZN(new_n470));
  INV_X1    g269(.A(new_n449), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n455), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n457), .B1(new_n473), .B2(new_n254), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n467), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n463), .A2(new_n471), .A3(new_n470), .A4(new_n468), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n444), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AND4_X1   g279(.A1(new_n444), .A2(new_n479), .A3(new_n475), .A4(new_n469), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n402), .B(new_n443), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n441), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n439), .A4(new_n440), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n442), .ZN(new_n486));
  INV_X1    g285(.A(new_n479), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n475), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n402), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n482), .A2(KEYINPUT92), .B1(KEYINPUT35), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT87), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n444), .A3(new_n479), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n402), .A4(new_n443), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT37), .B1(new_n472), .B2(new_n474), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n458), .A2(new_n498), .A3(new_n463), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n499), .A3(new_n467), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT38), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(KEYINPUT90), .A3(KEYINPUT38), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n441), .A2(new_n442), .A3(new_n477), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n453), .A2(new_n247), .A3(new_n455), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n446), .A2(new_n254), .A3(new_n448), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT37), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n499), .A3(new_n513), .A4(new_n467), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n419), .A2(new_n420), .ZN(new_n516));
  INV_X1    g315(.A(new_n408), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n424), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(new_n428), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT39), .B(new_n516), .C1(new_n520), .C2(new_n413), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n408), .B1(new_n429), .B2(new_n430), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n420), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n436), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT40), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n527), .A2(new_n528), .A3(new_n438), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n493), .A3(new_n492), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n283), .A2(new_n286), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n399), .A2(new_n401), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT36), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n283), .A2(KEYINPUT86), .A3(new_n286), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n486), .A2(new_n489), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n491), .A2(new_n496), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G43gat), .B(G50gat), .Z(new_n545));
  INV_X1    g344(.A(KEYINPUT15), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  NOR3_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n549), .B(new_n551), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(KEYINPUT94), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n552), .B2(KEYINPUT94), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n550), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(G1gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G1gat), .B2(new_n563), .ZN(new_n566));
  INV_X1    g365(.A(G8gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n571), .A2(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n562), .A2(KEYINPUT17), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(KEYINPUT18), .A3(new_n575), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n561), .B(new_n568), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n575), .B(KEYINPUT13), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT11), .B(G169gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n578), .A2(new_n592), .A3(new_n579), .A4(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n573), .A2(new_n571), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n561), .A2(new_n604), .B1(KEYINPUT41), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT101), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n613), .A2(new_n616), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G71gat), .B(G78gat), .Z(new_n621));
  XOR2_X1   g420(.A(KEYINPUT96), .B(G57gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G64gat), .ZN(new_n623));
  INV_X1    g422(.A(G64gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(G57gat), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT97), .Z(new_n628));
  INV_X1    g427(.A(new_n625), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n624), .A2(G57gat), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT9), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n626), .A2(new_n628), .B1(new_n621), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(KEYINPUT21), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT98), .ZN(new_n634));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n568), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT100), .Z(new_n640));
  XOR2_X1   g439(.A(new_n637), .B(new_n640), .Z(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n597), .A2(new_n603), .A3(new_n601), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n604), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n632), .A2(new_n604), .A3(KEYINPUT10), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n652), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  OAI211_X1 g465(.A(new_n663), .B(new_n666), .C1(new_n651), .C2(new_n656), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  INV_X1    g467(.A(new_n660), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n652), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n656), .A2(new_n651), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n620), .A2(new_n650), .A3(new_n674), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n544), .A2(new_n595), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n486), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(G1gat), .Z(G1324gat));
  INV_X1    g477(.A(new_n676), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n480), .A2(new_n481), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n567), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n676), .A2(new_n494), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n537), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n676), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n533), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n676), .B2(new_n690), .ZN(G1326gat));
  INV_X1    g490(.A(new_n541), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n402), .A2(new_n443), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT92), .B1(new_n680), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n496), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n532), .A2(new_n543), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n620), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n650), .A2(new_n595), .A3(new_n673), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n486), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT45), .Z(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n544), .B2(new_n620), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n700), .ZN(new_n708));
  INV_X1    g507(.A(new_n619), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n617), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n702), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n486), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n705), .A2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n703), .A2(G36gat), .A3(new_n494), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n713), .B2(new_n494), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1329gat));
  NOR3_X1   g518(.A1(new_n703), .A2(G43gat), .A3(new_n689), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT106), .ZN(new_n721));
  INV_X1    g520(.A(new_n537), .ZN(new_n722));
  OAI21_X1  g521(.A(G43gat), .B1(new_n713), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT47), .ZN(new_n724));
  OAI21_X1  g523(.A(G43gat), .B1(new_n713), .B2(new_n687), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g526(.A(G50gat), .B1(new_n713), .B2(new_n531), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n703), .A2(G50gat), .A3(new_n692), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n712), .A2(new_n541), .A3(new_n702), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n732), .B2(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g533(.A(new_n650), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n710), .A2(new_n594), .A3(new_n735), .A4(new_n674), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n708), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n486), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT107), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n622), .ZN(G1332gat));
  NOR2_X1   g541(.A1(new_n737), .A2(new_n494), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  NOR3_X1   g546(.A1(new_n737), .A2(G71gat), .A3(new_n689), .ZN(new_n748));
  INV_X1    g547(.A(new_n687), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(G71gat), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n738), .A2(new_n541), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n650), .A2(new_n594), .A3(new_n674), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n712), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n486), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n650), .A2(new_n594), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n701), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n673), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n739), .A2(new_n599), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  NOR3_X1   g563(.A1(new_n494), .A2(G92gat), .A3(new_n674), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n708), .A2(new_n710), .A3(new_n758), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n701), .B2(new_n758), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n712), .A2(new_n680), .A3(new_n755), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(new_n772), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT108), .B1(new_n773), .B2(G92gat), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(new_n761), .B2(new_n765), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n774), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n756), .B2(new_n687), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n689), .A2(G99gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n762), .B2(new_n783), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n674), .A2(G106gat), .A3(new_n531), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  INV_X1    g586(.A(new_n531), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n707), .A2(new_n788), .A3(new_n711), .A4(new_n755), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n707), .A2(new_n541), .A3(new_n711), .A4(new_n755), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n785), .B1(new_n767), .B2(new_n768), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n796), .B2(KEYINPUT53), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT111), .B(new_n787), .C1(new_n794), .C2(new_n795), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT112), .B(new_n791), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n669), .B2(new_n652), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n663), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n666), .B1(new_n670), .B2(new_n804), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n667), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n667), .C1(new_n808), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n808), .A2(new_n809), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n811), .A2(new_n594), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n580), .A2(new_n582), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT114), .Z(new_n817));
  NOR2_X1   g616(.A1(new_n574), .A2(new_n575), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n588), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n593), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n673), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n710), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n618), .B2(new_n619), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n735), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n675), .A2(new_n594), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n739), .A2(new_n829), .A3(new_n494), .A4(new_n402), .ZN(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n594), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n829), .B2(new_n692), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n834), .B(new_n541), .C1(new_n826), .C2(new_n828), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n680), .A2(new_n486), .A3(new_n689), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n594), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n838), .A2(KEYINPUT116), .A3(G113gat), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT116), .B1(new_n838), .B2(G113gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(G1340gat));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n837), .ZN(new_n842));
  OAI21_X1  g641(.A(G120gat), .B1(new_n842), .B2(new_n674), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n830), .A2(new_n293), .A3(new_n673), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  OAI21_X1  g644(.A(G127gat), .B1(new_n842), .B2(new_n735), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n289), .A3(new_n650), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n287), .A3(new_n710), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n710), .A3(new_n837), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n852), .A2(new_n853), .A3(G134gat), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n852), .B2(G134gat), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n850), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(new_n825), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n594), .A2(new_n814), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n821), .B1(new_n858), .B2(new_n810), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n620), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n620), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n857), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n827), .B1(new_n864), .B2(new_n735), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n865), .B2(new_n692), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n531), .B1(new_n826), .B2(new_n828), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n680), .A2(new_n537), .A3(new_n486), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n866), .A2(new_n594), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT119), .B1(new_n871), .B2(G141gat), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n749), .A2(new_n531), .A3(new_n680), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n829), .A2(new_n739), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(G141gat), .A3(new_n595), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n871), .B2(G141gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n872), .A2(new_n876), .A3(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  AOI221_X4 g677(.A(new_n875), .B1(KEYINPUT119), .B2(new_n878), .C1(new_n871), .C2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n874), .A2(new_n674), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n881), .A2(new_n882), .A3(G148gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n869), .A3(new_n870), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n674), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n650), .B1(new_n857), .B2(new_n860), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n868), .B(new_n541), .C1(new_n886), .C2(new_n827), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n867), .B2(new_n868), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n870), .A2(KEYINPUT59), .A3(new_n673), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n883), .B1(new_n890), .B2(G148gat), .ZN(G1345gat));
  INV_X1    g690(.A(new_n236), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n884), .B2(new_n735), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n735), .A2(new_n892), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n874), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n893), .B(new_n898), .C1(new_n874), .C2(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1346gat));
  NOR3_X1   g699(.A1(new_n874), .A2(G162gat), .A3(new_n620), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT121), .ZN(new_n902));
  OAI21_X1  g701(.A(G162gat), .B1(new_n884), .B2(new_n620), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n494), .A2(new_n739), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n689), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n836), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n595), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n905), .A2(new_n402), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n829), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(G169gat), .A3(new_n595), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT122), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n908), .B2(new_n674), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n674), .A2(G176gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n911), .B2(new_n916), .ZN(G1349gat));
  AND2_X1   g716(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n829), .A2(new_n345), .A3(new_n650), .A4(new_n910), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT123), .Z(new_n921));
  OAI211_X1 g720(.A(new_n650), .B(new_n907), .C1(new_n833), .C2(new_n835), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G183gat), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n918), .B(new_n919), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  AND4_X1   g723(.A1(KEYINPUT124), .A2(new_n921), .A3(KEYINPUT60), .A4(new_n923), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n836), .A2(new_n710), .A3(new_n907), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(G190gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n927), .B2(G190gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n710), .A2(new_n331), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n929), .A2(new_n930), .B1(new_n911), .B2(new_n931), .ZN(G1351gat));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(G197gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n749), .A2(new_n906), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n887), .B(new_n934), .C1(new_n867), .C2(new_n868), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n595), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n867), .A2(new_n934), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n595), .A2(new_n933), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1352gat));
  NOR3_X1   g738(.A1(new_n937), .A2(G204gat), .A3(new_n674), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n935), .B2(new_n674), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1353gat));
  INV_X1    g742(.A(new_n937), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n218), .A3(new_n650), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT126), .ZN(new_n946));
  OAI21_X1  g745(.A(G211gat), .B1(new_n935), .B2(new_n735), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT63), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT63), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G1354gat));
  AOI21_X1  g749(.A(G218gat), .B1(new_n944), .B2(new_n710), .ZN(new_n951));
  INV_X1    g750(.A(new_n935), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n710), .A2(G218gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(G1355gat));
endmodule


