//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G101), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n461), .A2(G137), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n461), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n460), .A2(new_n462), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n477), .B(new_n479), .C1(G124), .C2(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n482));
  OR2_X1    g057(.A1(G102), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n458), .B2(new_n459), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n459), .C2(new_n458), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G62), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(new_n498), .B1(G75), .B2(G543), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n496), .A2(KEYINPUT68), .A3(G62), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT5), .B(G543), .Z(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n501), .B2(KEYINPUT69), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n502), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n504), .A2(new_n505), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n503), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n496), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n524), .A2(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n496), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n495), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n527), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n496), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n495), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n516), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n503), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G651), .B1(new_n507), .B2(G91), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT71), .B(new_n551), .C1(new_n516), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n554), .B2(KEYINPUT9), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n509), .B(new_n555), .C1(new_n554), .C2(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(G299));
  INV_X1    g132(.A(G166), .ZN(G303));
  OR2_X1    g133(.A1(new_n496), .A2(G74), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n509), .B2(G49), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n507), .A2(new_n561), .A3(G87), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n561), .B1(new_n507), .B2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(G288));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n516), .B1(new_n525), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n496), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n495), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G305));
  INV_X1    g146(.A(G47), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT73), .B(G85), .Z(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n516), .B1(new_n525), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n496), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n495), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n574), .A2(KEYINPUT74), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  INV_X1    g155(.A(G54), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n516), .B2(KEYINPUT75), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n582), .B1(KEYINPUT75), .B2(new_n516), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT76), .B(G66), .Z(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n503), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n507), .A2(G92), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n583), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n580), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n580), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G286), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g171(.A(G299), .B(KEYINPUT77), .Z(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n595), .ZN(G297));
  AOI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n595), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g180(.A(KEYINPUT3), .B(G2104), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n463), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n461), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n480), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n462), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(G156));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT79), .Z(G401));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(G227));
  XOR2_X1   g222(.A(G1971), .B(G1976), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT19), .ZN(new_n649));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  AND2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT82), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n662), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n662), .B(new_n664), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(new_n666), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(G24), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G290), .B2(G16), .ZN(new_n675));
  INV_X1    g250(.A(G1986), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G25), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n461), .A2(G131), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n480), .A2(G119), .ZN(new_n681));
  OR2_X1    g256(.A1(G95), .A2(G2105), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n682), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n679), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT35), .B(G1991), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n675), .B2(new_n676), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n691));
  NAND2_X1  g266(.A1(G288), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g267(.A(KEYINPUT83), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n694), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n673), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n673), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1971), .ZN(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n570), .B2(G16), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT32), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1981), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n697), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n677), .B(new_n689), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT36), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n673), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n673), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT86), .Z(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT88), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n678), .A2(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n606), .A2(G127), .ZN(new_n721));
  NAND2_X1  g296(.A1(G115), .A2(G2104), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n462), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n720), .B(new_n723), .C1(G139), .C2(new_n461), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n678), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G2072), .Z(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G34), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n473), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n678), .A2(G27), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n678), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2078), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n733), .A2(G2084), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT89), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G301), .B2(new_n673), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G2078), .B2(new_n736), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT87), .B(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n748), .C1(new_n617), .C2(new_n678), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n732), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n726), .A2(new_n739), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n742), .A2(new_n743), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT90), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n717), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n678), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n480), .A2(G129), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT84), .Z(new_n758));
  AND2_X1   g333(.A1(new_n463), .A2(G105), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT26), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n759), .B(new_n761), .C1(G141), .C2(new_n461), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT85), .Z(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n678), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n716), .A2(new_n755), .A3(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT92), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n678), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n678), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT29), .Z(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n673), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n592), .B2(new_n673), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1348), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n673), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n541), .B2(new_n673), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1341), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n461), .A2(G140), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n480), .A2(G128), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n462), .A2(G116), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n678), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n774), .A2(new_n777), .A3(new_n780), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n673), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G1956), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n796), .B(new_n797), .C1(new_n772), .C2(new_n773), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n791), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n710), .A2(new_n769), .A3(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n804), .A2(new_n516), .B1(new_n525), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n496), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n495), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G860), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n592), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  INV_X1    g390(.A(new_n809), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n540), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n533), .B(new_n809), .C1(new_n538), .C2(new_n539), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT95), .Z(new_n823));
  OAI21_X1  g398(.A(new_n810), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n813), .B1(new_n823), .B2(new_n824), .ZN(G145));
  INV_X1    g400(.A(G37), .ZN(new_n826));
  XOR2_X1   g401(.A(G162), .B(new_n617), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n473), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n763), .A2(new_n724), .ZN(new_n829));
  INV_X1    g404(.A(new_n764), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n724), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n785), .B(G164), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n685), .ZN(new_n833));
  AOI22_X1  g408(.A1(G130), .A2(new_n480), .B1(new_n461), .B2(G142), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n837), .A2(new_n462), .A3(G118), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n462), .B2(G118), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n608), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n833), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n831), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n828), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT99), .B1(new_n845), .B2(new_n828), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n826), .B1(new_n828), .B2(new_n845), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(new_n816), .A2(new_n595), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n692), .A2(new_n693), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n570), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n577), .A2(KEYINPUT101), .A3(new_n578), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT101), .B1(new_n577), .B2(new_n578), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(G166), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n694), .A2(G305), .ZN(new_n859));
  OAI21_X1  g434(.A(G166), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n854), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n858), .A2(new_n860), .B1(new_n854), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT42), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n819), .B(new_n602), .Z(new_n865));
  AND2_X1   g440(.A1(new_n583), .A2(new_n587), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(G299), .C1(new_n590), .C2(new_n589), .ZN(new_n867));
  INV_X1    g442(.A(G299), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n591), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n591), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n864), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n852), .B1(new_n881), .B2(new_n595), .ZN(G295));
  OAI21_X1  g457(.A(new_n852), .B1(new_n881), .B2(new_n595), .ZN(G331));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n817), .A2(new_n818), .A3(G301), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G301), .B1(new_n817), .B2(new_n818), .ZN(new_n887));
  OAI21_X1  g462(.A(G286), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(G168), .A3(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n871), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n888), .B(new_n890), .C1(new_n874), .C2(new_n878), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n863), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n863), .A2(new_n892), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n826), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n902), .A2(new_n890), .A3(new_n888), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n870), .B1(new_n891), .B2(new_n873), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n863), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n900), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n884), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT102), .B1(new_n898), .B2(KEYINPUT43), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(KEYINPUT44), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n900), .A2(new_n907), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n896), .A2(new_n908), .A3(new_n826), .A4(new_n897), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  AOI22_X1  g491(.A1(KEYINPUT43), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n912), .A2(new_n919), .ZN(G397));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  INV_X1    g496(.A(new_n493), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n492), .B1(new_n606), .B2(new_n489), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n924), .B2(new_n487), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n468), .A2(new_n472), .A3(G40), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n763), .A3(G1996), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT106), .Z(new_n931));
  XOR2_X1   g506(.A(new_n785), .B(G2067), .Z(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n830), .B2(G1996), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n933), .B2(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n684), .B(new_n687), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT105), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n921), .C1(new_n924), .C2(new_n487), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(KEYINPUT108), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n925), .A2(new_n947), .A3(KEYINPUT50), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n468), .A2(new_n472), .A3(G40), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n750), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n928), .B1(new_n925), .B2(new_n926), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n925), .A2(new_n926), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n714), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n950), .B1(new_n949), .B2(new_n953), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT122), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G286), .A2(G8), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT123), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n949), .A2(new_n953), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT115), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT122), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n958), .A4(new_n954), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n959), .A2(new_n960), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT125), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT125), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n974), .B(G8), .C1(new_n959), .C2(new_n960), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n972), .A2(new_n973), .A3(new_n963), .A4(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n961), .A2(G8), .A3(new_n968), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n977), .B2(new_n963), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(KEYINPUT124), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT124), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(new_n973), .C1(new_n977), .C2(new_n963), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n969), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT62), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n969), .C1(new_n979), .C2(new_n981), .ZN(new_n985));
  NOR2_X1   g560(.A1(G164), .A2(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n951), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n694), .B2(G1976), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  NAND2_X1  g567(.A1(G288), .A2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n988), .B(new_n993), .C1(new_n694), .C2(G1976), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n994), .B2(KEYINPUT52), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n570), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT49), .B1(new_n996), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(new_n988), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n989), .A2(new_n990), .A3(new_n1005), .A4(new_n993), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n995), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1008));
  NAND3_X1  g583(.A1(G303), .A2(G8), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(G166), .B2(new_n971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT107), .B1(new_n925), .B2(new_n926), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n986), .A2(new_n1014), .A3(KEYINPUT45), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n955), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1971), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n949), .A2(new_n951), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(G2090), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n943), .A2(new_n951), .A3(new_n945), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(G2090), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n971), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1012), .A2(new_n1024), .A3(KEYINPUT114), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1024), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1007), .A2(new_n1021), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1019), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n949), .A2(KEYINPUT118), .A3(new_n951), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n743), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1016), .A2(G2078), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1032), .A2(KEYINPUT53), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n956), .A2(new_n957), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT53), .A3(new_n738), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1027), .A2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n983), .A2(new_n985), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n987), .A2(G2067), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT118), .B1(new_n949), .B2(new_n951), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1028), .B(new_n928), .C1(new_n946), .C2(new_n948), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1348), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT121), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1029), .A2(new_n1045), .A3(new_n1030), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1041), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(KEYINPUT121), .A3(new_n1050), .A4(new_n1047), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1040), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT60), .A3(new_n592), .A4(new_n1051), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1013), .A2(new_n955), .A3(new_n1015), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1022), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT117), .B1(new_n1022), .B2(new_n1061), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1060), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(G299), .B(KEYINPUT57), .Z(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1067), .B(new_n1060), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1058), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n987), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1016), .B2(G1996), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n540), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1076), .B(new_n1077), .C1(KEYINPUT119), .C2(KEYINPUT59), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1053), .A2(new_n1057), .A3(new_n1073), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1069), .B1(new_n1046), .B2(new_n591), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1070), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1032), .A2(KEYINPUT53), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1031), .A2(new_n1033), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n1089), .B2(G301), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1036), .A2(G171), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1031), .A2(new_n1033), .A3(G301), .A4(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT54), .B1(new_n1037), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1092), .A2(new_n1027), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1087), .A2(new_n1095), .A3(new_n982), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n988), .B(KEYINPUT112), .Z(new_n1097));
  NOR2_X1   g672(.A1(G288), .A2(G1976), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT113), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1100));
  INV_X1    g675(.A(new_n998), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1007), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1021), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1007), .A2(new_n1021), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1020), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1012), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n970), .A2(new_n971), .A3(G286), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1105), .A2(new_n1109), .A3(KEYINPUT63), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1110), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1027), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1104), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1096), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n942), .B1(new_n1039), .B2(new_n1116), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n935), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT46), .B1(new_n935), .B2(G1996), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n932), .A2(new_n758), .A3(new_n762), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1118), .A2(new_n1119), .B1(new_n929), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT47), .Z(new_n1122));
  NOR2_X1   g697(.A1(new_n785), .A2(G2067), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n685), .A2(new_n687), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT126), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n934), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1122), .B1(new_n1126), .B2(new_n935), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n937), .B(KEYINPUT127), .Z(new_n1128));
  NOR2_X1   g703(.A1(new_n939), .A2(new_n935), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1117), .A2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g707(.A(new_n634), .ZN(new_n1134));
  INV_X1    g708(.A(G319), .ZN(new_n1135));
  NOR3_X1   g709(.A1(new_n1134), .A2(new_n1135), .A3(G227), .ZN(new_n1136));
  AND3_X1   g710(.A1(new_n668), .A2(new_n670), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g711(.A(new_n1137), .B(new_n850), .C1(new_n910), .C2(new_n911), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


