//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g0003(.A(KEYINPUT64), .B1(new_n203), .B2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n206), .A2(new_n207), .A3(new_n201), .A4(new_n202), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n212), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT66), .B(G244), .Z(new_n225));
  AND2_X1   g0025(.A1(new_n225), .A2(G77), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n217), .B(new_n224), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n207), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n245), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(KEYINPUT81), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n256), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  INV_X1    g0063(.A(G87), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n262), .A2(new_n263), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G226), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n255), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT67), .A2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT67), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n222), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n253), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n280), .B2(new_n275), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n255), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n276), .A2(new_n279), .B1(new_n282), .B2(G232), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n270), .A2(G179), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n270), .B2(new_n283), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n222), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n266), .B2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n258), .A2(new_n260), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n202), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G58), .A2(G68), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT76), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n203), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(G159), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n290), .B1(new_n306), .B2(KEYINPUT16), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT78), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT78), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n258), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n260), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n291), .A2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT77), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n257), .A2(G33), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n212), .B1(new_n308), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n317), .B2(new_n291), .ZN(new_n318));
  AOI21_X1  g0118(.A(G20), .B1(new_n258), .B2(new_n260), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n319), .A2(KEYINPUT77), .A3(KEYINPUT7), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n314), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n305), .B1(new_n321), .B2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n307), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT8), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n201), .B2(KEYINPUT70), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT8), .A3(G58), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n211), .A2(G20), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT79), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n222), .A3(new_n288), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n330), .B2(KEYINPUT79), .ZN(new_n334));
  INV_X1    g0134(.A(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(new_n328), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n331), .A2(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n287), .B1(new_n323), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n252), .B1(new_n338), .B2(KEYINPUT18), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n270), .A2(G179), .A3(new_n283), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n270), .A2(new_n283), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n285), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n319), .A2(KEYINPUT7), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n291), .B(G20), .C1(new_n258), .C2(new_n260), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n303), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n289), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT77), .B1(new_n319), .B2(KEYINPUT7), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n315), .B(new_n291), .C1(new_n266), .C2(G20), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n312), .B2(new_n313), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n202), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n348), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n337), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT18), .B(new_n342), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT80), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n338), .A2(new_n358), .A3(KEYINPUT18), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n349), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(new_n307), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT81), .B(new_n360), .C1(new_n362), .C2(new_n287), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n339), .A2(new_n357), .A3(new_n359), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n270), .B2(new_n283), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G190), .B2(new_n341), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT17), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n276), .A2(new_n279), .B1(new_n282), .B2(G226), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n267), .A2(new_n263), .B1(new_n205), .B2(new_n266), .ZN(new_n372));
  INV_X1    g0172(.A(G222), .ZN(new_n373));
  OR3_X1    g0173(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT69), .B1(new_n262), .B2(new_n373), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n376), .B2(new_n254), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n212), .A2(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT71), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(KEYINPUT71), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n328), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G150), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n304), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n212), .B1(new_n204), .B2(new_n208), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n289), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n333), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n207), .B1(new_n211), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n388), .A2(new_n389), .B1(new_n207), .B2(new_n335), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT9), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(KEYINPUT9), .A3(new_n390), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n379), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n378), .A2(new_n365), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT10), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n392), .A2(new_n393), .ZN(new_n397));
  INV_X1    g0197(.A(new_n395), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT10), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n379), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n276), .A2(new_n279), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n282), .A2(new_n225), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G107), .ZN(new_n407));
  INV_X1    g0207(.A(G232), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n406), .B1(new_n407), .B2(new_n266), .C1(new_n408), .C2(new_n262), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n255), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n411), .B2(G179), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(KEYINPUT73), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n329), .A2(G77), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n333), .A2(new_n416), .B1(G77), .B2(new_n332), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G20), .A2(G77), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT8), .B(G58), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n418), .B1(new_n419), .B2(new_n380), .C1(new_n304), .C2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n289), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n411), .B2(new_n285), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n410), .B2(new_n365), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT72), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n410), .B2(G190), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n410), .A2(new_n425), .A3(G190), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n415), .A2(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n377), .A2(new_n285), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n387), .A2(new_n390), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(G179), .C2(new_n377), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n401), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n382), .A2(G77), .A3(new_n381), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n303), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n290), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(KEYINPUT11), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n329), .A2(G68), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n333), .B2(new_n439), .ZN(new_n440));
  OR3_X1    g0240(.A1(new_n333), .A2(new_n438), .A3(new_n439), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n436), .A2(KEYINPUT11), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n335), .A2(new_n202), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT12), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT75), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G97), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n262), .B2(new_n268), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n267), .A2(new_n408), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n255), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n276), .A2(new_n279), .B1(new_n282), .B2(G238), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT14), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(G169), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n413), .B2(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n458), .B2(G169), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n447), .B(new_n448), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n447), .A2(new_n448), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(G200), .ZN(new_n465));
  INV_X1    g0265(.A(G190), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n458), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n370), .A2(new_n433), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(new_n266), .A3(KEYINPUT4), .A4(G244), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AND4_X1   g0277(.A1(new_n258), .A2(new_n256), .A3(new_n260), .A4(new_n261), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT4), .B1(new_n478), .B2(G244), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n255), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n272), .B2(new_n273), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n211), .B(G45), .C1(new_n481), .C2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n255), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT67), .A2(G41), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT5), .B1(new_n486), .B2(new_n271), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n483), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n485), .A2(G257), .B1(new_n488), .B2(new_n279), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n285), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n480), .A2(new_n413), .A3(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n321), .A2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n407), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n407), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G20), .B1(G77), .B2(new_n303), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n290), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n335), .A2(new_n495), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n388), .B1(G1), .B2(new_n259), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n495), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n491), .B(new_n492), .C1(new_n501), .C2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n258), .A2(new_n260), .A3(new_n212), .A4(G87), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n266), .A2(new_n212), .A3(new_n508), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n212), .B2(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n407), .A2(KEYINPUT23), .A3(G20), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n512), .A2(new_n521), .A3(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n289), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n333), .B1(new_n211), .B2(G33), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n332), .B2(G107), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n332), .A2(new_n526), .A3(G107), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n525), .A2(G107), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n258), .A2(new_n260), .A3(G257), .A4(G1698), .ZN(new_n531));
  INV_X1    g0331(.A(G294), .ZN(new_n532));
  INV_X1    g0332(.A(G250), .ZN(new_n533));
  OAI221_X1 g0333(.A(new_n531), .B1(new_n259), .B2(new_n532), .C1(new_n262), .C2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n255), .B1(G264), .B2(new_n485), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n482), .A2(new_n279), .A3(new_n484), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(G190), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n531), .B1(new_n259), .B2(new_n532), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n262), .A2(new_n533), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n255), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n485), .A2(G264), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n524), .A2(new_n530), .A3(new_n537), .A4(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n500), .B1(new_n352), .B2(new_n407), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n504), .B1(new_n545), .B2(new_n289), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n480), .A2(new_n466), .A3(new_n489), .ZN(new_n547));
  AOI21_X1  g0347(.A(G200), .B1(new_n480), .B2(new_n489), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n505), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n332), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n525), .B2(new_n552), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n288), .A2(new_n222), .B1(G20), .B2(new_n552), .ZN(new_n555));
  AOI21_X1  g0355(.A(G20), .B1(G33), .B2(G283), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n259), .A2(G97), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT86), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT86), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT20), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT86), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT20), .B1(new_n566), .B2(new_n555), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n554), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G169), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n258), .A2(new_n260), .A3(G257), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n473), .B1(G303), .B2(new_n293), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n266), .A2(G264), .A3(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n254), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G270), .B(new_n254), .C1(new_n487), .C2(new_n483), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n536), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n536), .A3(KEYINPUT85), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n551), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n568), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n266), .A2(G257), .ZN(new_n582));
  INV_X1    g0382(.A(new_n473), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n266), .ZN(new_n585));
  INV_X1    g0385(.A(new_n572), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n255), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n574), .A2(new_n536), .A3(KEYINPUT85), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT85), .B1(new_n574), .B2(new_n536), .ZN(new_n589));
  OAI211_X1 g0389(.A(G190), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n581), .B(new_n590), .C1(new_n579), .C2(new_n365), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(KEYINPUT21), .A3(G169), .A4(new_n568), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n579), .A2(G179), .A3(new_n568), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n580), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n503), .A2(new_n419), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n419), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n332), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n258), .A2(new_n260), .A3(new_n212), .A4(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n380), .B2(new_n495), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n212), .B1(new_n449), .B2(new_n602), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n497), .A2(new_n264), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT83), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n289), .B1(new_n610), .B2(KEYINPUT84), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n606), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n601), .B(new_n603), .C1(new_n612), .C2(new_n607), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT84), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n597), .B(new_n600), .C1(new_n611), .C2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n473), .A2(new_n266), .A3(G238), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(G1698), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n513), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n255), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n275), .A2(G1), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n254), .A2(G274), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n533), .B1(new_n211), .B2(G45), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n254), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT82), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n254), .A3(KEYINPUT82), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n620), .A2(new_n413), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n618), .A2(new_n513), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n473), .A2(new_n266), .A3(G238), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n254), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n622), .ZN(new_n633));
  INV_X1    g0433(.A(new_n627), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT82), .B1(new_n623), .B2(new_n254), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n285), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n616), .A2(new_n629), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n542), .A2(new_n285), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n535), .A2(new_n413), .A3(new_n536), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n290), .B1(new_n520), .B2(new_n522), .ZN(new_n641));
  INV_X1    g0441(.A(new_n530), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n620), .A2(new_n466), .A3(new_n628), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n632), .A2(new_n636), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(G200), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n290), .B1(new_n613), .B2(new_n614), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n610), .A2(KEYINPUT84), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n599), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n525), .A2(G87), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n638), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n550), .A2(new_n595), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n470), .A2(new_n653), .ZN(G372));
  INV_X1    g0454(.A(KEYINPUT17), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n368), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n415), .A2(new_n423), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n467), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n656), .B1(new_n463), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n342), .B1(new_n354), .B2(new_n355), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n360), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n356), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n401), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n432), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n637), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n620), .A2(new_n628), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .A3(new_n285), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n668), .B1(new_n673), .B2(new_n629), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT88), .B1(new_n671), .B2(new_n285), .ZN(new_n675));
  AOI211_X1 g0475(.A(new_n669), .B(G169), .C1(new_n620), .C2(new_n628), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n668), .B(new_n629), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n616), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n505), .A2(new_n544), .A3(new_n549), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT90), .A4(new_n651), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n643), .A2(new_n580), .A3(new_n593), .A4(new_n594), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n651), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n629), .B1(new_n675), .B2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n677), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n687), .B2(new_n616), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT90), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n596), .B(new_n599), .C1(new_n647), .C2(new_n648), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n637), .A2(new_n629), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n600), .B(new_n650), .C1(new_n611), .C2(new_n615), .ZN(new_n693));
  AOI21_X1  g0493(.A(G200), .B1(new_n620), .B2(new_n628), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n466), .B2(new_n645), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n691), .A2(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n696), .B2(new_n505), .ZN(new_n697));
  INV_X1    g0497(.A(new_n505), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n679), .B(new_n697), .C1(new_n699), .C2(KEYINPUT26), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n667), .B1(new_n469), .B2(new_n701), .ZN(G369));
  NAND3_X1  g0502(.A1(new_n580), .A2(new_n593), .A3(new_n594), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n581), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n595), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n643), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n709), .B1(new_n641), .B2(new_n642), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n544), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n643), .A2(new_n709), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n703), .A2(new_n710), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n718), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n215), .ZN(new_n727));
  INV_X1    g0527(.A(new_n274), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n606), .A2(G116), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n220), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT26), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n696), .B2(new_n505), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT94), .B(new_n735), .C1(new_n696), .C2(new_n505), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n691), .B1(new_n686), .B2(new_n677), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n741), .A2(new_n735), .A3(new_n505), .A4(new_n684), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n505), .A2(new_n744), .A3(new_n549), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(new_n505), .B2(new_n549), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n544), .B(new_n682), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n679), .B1(new_n747), .B2(new_n684), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n710), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(new_n710), .C1(new_n690), .C2(new_n700), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n671), .A2(new_n413), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n579), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n592), .A2(KEYINPUT93), .A3(new_n413), .A4(new_n671), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(new_n490), .A4(new_n542), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n540), .A2(new_n541), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT91), .B1(new_n759), .B2(new_n671), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT91), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n645), .A2(new_n761), .A3(new_n535), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(G179), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n490), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT92), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(KEYINPUT92), .B(KEYINPUT30), .C1(new_n763), .C2(new_n765), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n709), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(new_n653), .B2(new_n710), .ZN(new_n772));
  OAI211_X1 g0572(.A(KEYINPUT31), .B(new_n709), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n753), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n734), .B1(new_n777), .B2(G1), .ZN(G364));
  AND2_X1   g0578(.A1(new_n212), .A2(G13), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n211), .B1(new_n779), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n729), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n713), .A2(G330), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n714), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT97), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n785), .B1(new_n787), .B2(G20), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n786), .A2(KEYINPUT97), .A3(new_n212), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n222), .B1(G20), .B2(new_n285), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n727), .A2(new_n266), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G45), .B2(new_n220), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n275), .C2(new_n250), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n727), .A2(new_n293), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n552), .B2(new_n727), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n793), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G179), .A2(G200), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n212), .B1(new_n802), .B2(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n532), .ZN(new_n804));
  NAND3_X1  g0604(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G190), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(KEYINPUT33), .A2(G317), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(KEYINPUT33), .A2(G317), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n805), .A2(new_n466), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n804), .B(new_n811), .C1(G326), .C2(new_n812), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n212), .A2(KEYINPUT98), .A3(G190), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT98), .B1(new_n212), .B2(G190), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G329), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n212), .A2(new_n466), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n413), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n293), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n365), .A2(G179), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n212), .A2(G190), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n820), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n825), .A2(new_n584), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n814), .A2(new_n815), .A3(new_n824), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n823), .B(new_n829), .C1(G283), .C2(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n813), .A2(new_n818), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n830), .A2(new_n407), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n201), .A2(new_n821), .B1(new_n825), .B2(new_n264), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n266), .B1(new_n827), .B2(new_n205), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n812), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n807), .A2(new_n202), .B1(new_n840), .B2(new_n207), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n803), .A2(new_n495), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT32), .B1(new_n816), .B2(new_n302), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n816), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n839), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n835), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n801), .B1(new_n848), .B2(new_n791), .ZN(new_n849));
  INV_X1    g0649(.A(new_n790), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n713), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n784), .B1(new_n851), .B2(new_n782), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n853));
  XNOR2_X1  g0653(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  OR2_X1    g0655(.A1(new_n710), .A2(new_n422), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n657), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n429), .A2(new_n856), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n701), .B2(new_n709), .ZN(new_n860));
  INV_X1    g0660(.A(new_n859), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n710), .B(new_n861), .C1(new_n690), .C2(new_n700), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n782), .B1(new_n863), .B2(new_n775), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n775), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n791), .A2(new_n786), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n782), .B1(G77), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n821), .ZN(new_n869));
  INV_X1    g0669(.A(new_n827), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G143), .A2(new_n869), .B1(new_n870), .B2(G159), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n871), .B1(new_n840), .B2(new_n872), .C1(new_n384), .C2(new_n807), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT34), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n831), .A2(G68), .ZN(new_n877));
  INV_X1    g0677(.A(new_n825), .ZN(new_n878));
  INV_X1    g0678(.A(new_n803), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(G50), .B1(new_n879), .B2(G58), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(G132), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n266), .B1(new_n816), .B2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT103), .Z(new_n884));
  AOI21_X1  g0684(.A(new_n842), .B1(new_n812), .B2(G303), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT102), .B(G283), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n807), .B2(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n821), .A2(new_n532), .B1(new_n827), .B2(new_n552), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n266), .B(new_n888), .C1(G107), .C2(new_n878), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n831), .A2(G87), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n889), .B(new_n890), .C1(new_n828), .C2(new_n816), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n881), .A2(new_n884), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n868), .B1(new_n892), .B2(new_n791), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n861), .B2(new_n787), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n865), .A2(new_n894), .ZN(G384));
  OR2_X1    g0695(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n223), .A4(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  NAND4_X1  g0699(.A1(new_n221), .A2(G77), .A3(new_n298), .A4(new_n299), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n211), .B(G13), .C1(new_n900), .C2(new_n246), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n666), .B1(new_n753), .B2(new_n470), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT106), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n349), .B1(new_n306), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n295), .A2(new_n305), .A3(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n307), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n337), .ZN(new_n910));
  INV_X1    g0710(.A(new_n707), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n364), .B2(new_n369), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n910), .A2(new_n342), .B1(new_n362), .B2(new_n367), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n912), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n354), .B2(new_n355), .ZN(new_n917));
  AND4_X1   g0717(.A1(new_n914), .A2(new_n368), .A3(new_n661), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n913), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n664), .B2(new_n656), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n661), .A2(new_n368), .A3(new_n917), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT37), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n905), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n916), .A2(new_n918), .ZN(new_n928));
  OAI211_X1 g0728(.A(KEYINPUT38), .B(new_n928), .C1(new_n370), .C2(new_n912), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n913), .B2(new_n919), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n463), .A2(new_n709), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n447), .A2(new_n448), .A3(new_n709), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT104), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n468), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n658), .A2(new_n710), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n862), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n929), .A2(new_n930), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n664), .A2(new_n707), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n904), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n921), .A2(new_n926), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n859), .B1(new_n772), .B2(new_n773), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n463), .A2(new_n467), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(new_n938), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT40), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n942), .A2(new_n953), .A3(new_n950), .A4(new_n948), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n470), .A3(new_n774), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n470), .A2(new_n774), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n952), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(G330), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n211), .B2(new_n779), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n946), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n902), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NOR3_X1   g0763(.A1(new_n241), .A2(new_n727), .A3(new_n266), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n792), .B1(new_n215), .B2(new_n419), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n782), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G150), .A2(new_n869), .B1(new_n870), .B2(G50), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n266), .C1(new_n201), .C2(new_n825), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n803), .A2(new_n202), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(G143), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n970), .B1(new_n840), .B2(new_n971), .C1(new_n302), .C2(new_n807), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n830), .A2(new_n205), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n816), .A2(new_n872), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n968), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT109), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n825), .A2(new_n552), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n977), .A2(KEYINPUT46), .B1(new_n532), .B2(new_n807), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G311), .B2(new_n812), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n827), .A2(new_n886), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n266), .B(new_n980), .C1(G303), .C2(new_n869), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n977), .A2(KEYINPUT46), .B1(G107), .B2(new_n879), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT108), .B(G317), .Z(new_n983));
  AOI22_X1  g0783(.A1(G97), .A2(new_n831), .B1(new_n817), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n966), .B1(new_n987), .B2(new_n791), .ZN(new_n988));
  INV_X1    g0788(.A(new_n693), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n688), .B1(new_n989), .B2(new_n710), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n741), .A2(new_n693), .A3(new_n709), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n850), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n546), .A2(new_n710), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n505), .A2(new_n549), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT95), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n505), .A2(new_n549), .A3(new_n744), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n698), .B2(new_n709), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n719), .A2(new_n724), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n999), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n505), .B1(new_n1005), .B2(new_n643), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1003), .A2(KEYINPUT42), .B1(new_n710), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT107), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT107), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1004), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n992), .B(KEYINPUT43), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n1012), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n722), .A2(new_n1000), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n725), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n1000), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT45), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1000), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n721), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n722), .A3(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n719), .B(new_n723), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(new_n714), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n777), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1033), .A2(new_n776), .A3(new_n753), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n729), .B(KEYINPUT41), .Z(new_n1035));
  OAI21_X1  g0835(.A(new_n780), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n994), .B1(new_n1019), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(G387));
  NAND2_X1  g0838(.A1(new_n1031), .A2(new_n781), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n782), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n731), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n799), .A2(new_n1041), .B1(new_n407), .B2(new_n727), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n238), .A2(new_n275), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n420), .A2(G50), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT50), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n731), .B(new_n275), .C1(new_n202), .C2(new_n205), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n794), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1042), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1040), .B1(new_n1048), .B2(new_n792), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n879), .A2(new_n598), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n840), .B2(new_n302), .C1(new_n336), .C2(new_n807), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G50), .A2(new_n869), .B1(new_n870), .B2(G68), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n293), .B1(new_n878), .B2(G77), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n495), .C2(new_n830), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(G150), .C2(new_n817), .ZN(new_n1055));
  INV_X1    g0855(.A(G326), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n293), .B1(new_n816), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n869), .A2(new_n983), .B1(new_n870), .B2(G303), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n840), .B2(new_n822), .C1(new_n828), .C2(new_n807), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n825), .A2(new_n532), .B1(new_n803), .B2(new_n886), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT110), .Z(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1057), .B(new_n1067), .C1(G116), .C2(new_n831), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1055), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n791), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1049), .B1(new_n719), .B2(new_n850), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1032), .A2(new_n729), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n777), .A2(new_n1031), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1039), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(G393));
  AND2_X1   g0875(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1076), .A2(new_n1033), .A3(new_n730), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1027), .A2(new_n781), .A3(new_n1028), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1000), .A2(new_n790), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n793), .B1(G97), .B2(new_n727), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n794), .A2(new_n245), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1040), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n879), .A2(G116), .B1(G303), .B2(new_n806), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT111), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n816), .A2(new_n822), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n293), .B1(new_n827), .B2(new_n532), .C1(new_n825), .C2(new_n886), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1084), .A2(new_n836), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n869), .A2(G311), .B1(G317), .B2(new_n812), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT52), .Z(new_n1089));
  OAI21_X1  g0889(.A(new_n890), .B1(new_n971), .B2(new_n816), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n266), .B1(new_n827), .B2(new_n420), .C1(new_n202), .C2(new_n825), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n807), .A2(new_n207), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n803), .A2(new_n205), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n840), .A2(new_n384), .B1(new_n821), .B2(new_n302), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1087), .A2(new_n1089), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1079), .B(new_n1082), .C1(new_n1071), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT112), .B1(new_n1078), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1078), .A2(KEYINPUT112), .A3(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1077), .B1(new_n1099), .B2(new_n1100), .ZN(G390));
  NOR2_X1   g0901(.A1(new_n775), .A2(new_n469), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT114), .B1(new_n903), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n469), .B1(new_n750), .B2(new_n752), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT114), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1105), .A2(new_n1102), .A3(new_n1106), .A4(new_n666), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n774), .A2(G330), .A3(new_n861), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n939), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n948), .A2(new_n950), .A3(G330), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n862), .A2(new_n940), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT115), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n940), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n738), .B(new_n739), .C1(new_n699), .C2(new_n735), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n682), .A2(new_n544), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n997), .B2(new_n998), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n741), .B1(new_n1119), .B2(new_n651), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n709), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1116), .B1(new_n1121), .B2(new_n861), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT115), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n948), .A2(new_n950), .A3(G330), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n950), .B1(new_n948), .B2(G330), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n1113), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1115), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1111), .A2(KEYINPUT113), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n932), .B1(new_n941), .B2(new_n935), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n947), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1131), .B(new_n934), .C1(new_n1122), .C2(new_n939), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1130), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1108), .B(new_n1128), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1133), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n679), .A2(new_n680), .A3(new_n651), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT90), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n682), .A3(new_n681), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n697), .A2(new_n679), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n741), .A2(new_n505), .A3(new_n684), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n735), .ZN(new_n1143));
  AOI211_X1 g0943(.A(KEYINPUT29), .B(new_n709), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n997), .A2(new_n998), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n688), .A3(new_n544), .A4(new_n682), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n679), .C1(new_n742), .C2(new_n740), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n751), .B1(new_n1147), .B2(new_n710), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n470), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n1103), .A3(new_n667), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1106), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n903), .A2(KEYINPUT114), .A3(new_n1103), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1127), .A2(new_n1123), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1124), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1151), .B(new_n1152), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1136), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1135), .A2(new_n1156), .A3(new_n729), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n781), .B1(new_n1134), .B2(new_n1133), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n782), .B1(new_n328), .B2(new_n867), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n266), .B1(new_n827), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n878), .A2(G150), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1163));
  OAI22_X1  g0963(.A1(new_n1162), .A2(new_n1163), .B1(new_n872), .B2(new_n807), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(G132), .C2(new_n869), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n879), .A2(G159), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1162), .A2(new_n1163), .B1(new_n812), .B2(G128), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G50), .A2(new_n831), .B1(new_n817), .B2(G125), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT117), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n821), .A2(new_n552), .B1(new_n827), .B2(new_n495), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n266), .B(new_n1171), .C1(G87), .C2(new_n878), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n807), .A2(new_n407), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1093), .B(new_n1173), .C1(G283), .C2(new_n812), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n817), .A2(G294), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n877), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1169), .A2(KEYINPUT117), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1170), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1159), .B1(new_n1178), .B2(new_n791), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n932), .B2(new_n786), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT118), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1158), .A2(KEYINPUT119), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT119), .B1(new_n1158), .B2(new_n1183), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1157), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1157), .B(KEYINPUT120), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(G378));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n936), .A2(new_n943), .A3(new_n944), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n401), .A2(new_n432), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n707), .B1(new_n387), .B2(new_n390), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR3_X1    g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n955), .B2(G330), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n955), .A2(G330), .A3(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1192), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1205), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n945), .B1(new_n1207), .B2(new_n1203), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1191), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT122), .B1(new_n1135), .B2(new_n1108), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT122), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1129), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1130), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1211), .B(new_n1212), .C1(new_n1217), .C2(new_n1128), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1209), .B1(new_n1210), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1108), .B1(new_n1136), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1211), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1135), .A2(KEYINPUT122), .A3(new_n1108), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1219), .B(new_n729), .C1(new_n1225), .C2(KEYINPUT57), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1200), .A2(new_n786), .A3(new_n1201), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n782), .B1(G50), .B2(new_n867), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n274), .B2(new_n293), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n970), .B1(new_n807), .B2(new_n495), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n274), .B(new_n293), .C1(new_n821), .C2(new_n407), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n825), .A2(new_n205), .B1(new_n827), .B2(new_n419), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G283), .C2(new_n817), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n831), .A2(G58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1231), .B(new_n1236), .C1(G116), .C2(new_n812), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1230), .B1(new_n1237), .B2(KEYINPUT58), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n807), .A2(new_n882), .B1(new_n803), .B2(new_n384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n870), .A2(G137), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n821), .C1(new_n825), .C2(new_n1160), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1239), .B(new_n1242), .C1(G125), .C2(new_n812), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n259), .B(new_n280), .C1(new_n830), .C2(new_n302), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G124), .B2(new_n817), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT59), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1238), .B1(KEYINPUT58), .B2(new_n1237), .C1(new_n1245), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1228), .B1(new_n1250), .B2(new_n791), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1227), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1220), .B2(new_n780), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT121), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT121), .B(new_n1252), .C1(new_n1220), .C2(new_n780), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1226), .A2(new_n1257), .ZN(G375));
  XNOR2_X1  g1058(.A(new_n780), .B(KEYINPUT123), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1221), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1040), .B1(new_n202), .B2(new_n866), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G283), .A2(new_n869), .B1(new_n870), .B2(G107), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n293), .C1(new_n495), .C2(new_n825), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n973), .B(new_n1263), .C1(G303), .C2(new_n817), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1050), .B1(new_n840), .B2(new_n532), .C1(new_n552), .C2(new_n807), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n812), .A2(G132), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT124), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1235), .B1(new_n1241), .B2(new_n816), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n807), .A2(new_n1160), .B1(new_n803), .B2(new_n207), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n266), .B1(new_n827), .B2(new_n384), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n872), .A2(new_n821), .B1(new_n825), .B2(new_n302), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1264), .A2(new_n1266), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1261), .B1(new_n1274), .B2(new_n1071), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n939), .B2(new_n786), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1260), .A2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1035), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1155), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1278), .B2(new_n1280), .ZN(G381));
  OR2_X1    g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  OR4_X1    g1082(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G381), .ZN(new_n1284));
  INV_X1    g1084(.A(G375), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1157), .A2(new_n1183), .A3(new_n1158), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n708), .A2(G213), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1285), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(new_n1290), .A3(G213), .ZN(G409));
  NAND3_X1  g1091(.A1(G378), .A2(new_n1226), .A3(new_n1257), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1279), .B1(new_n1210), .B2(new_n1218), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1220), .B1(new_n1293), .B2(new_n1259), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1252), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1286), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1288), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1278), .B1(KEYINPUT60), .B2(new_n1155), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1212), .A2(new_n1221), .A3(KEYINPUT60), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n729), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1277), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G384), .B(KEYINPUT125), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  OAI221_X1 g1104(.A(new_n1277), .B1(KEYINPUT125), .B2(G384), .C1(new_n1299), .C2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G2897), .A3(new_n1289), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1289), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1289), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1306), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1297), .A2(new_n1288), .A3(new_n1315), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1312), .A2(new_n1316), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1282), .ZN(new_n1320));
  AND2_X1   g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(G390), .ZN(new_n1323));
  OAI221_X1 g1123(.A(new_n1077), .B1(new_n1099), .B2(new_n1100), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1037), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1037), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1330), .B(new_n1327), .C1(new_n1313), .C2(new_n1310), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1289), .B(new_n1306), .C1(new_n1292), .C2(new_n1296), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT126), .B1(new_n1333), .B2(KEYINPUT63), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(KEYINPUT63), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1317), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1332), .A2(new_n1334), .A3(new_n1335), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1329), .A2(new_n1339), .ZN(G405));
  NAND2_X1  g1140(.A1(G375), .A2(new_n1286), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1292), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1315), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1292), .A3(new_n1306), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1346), .B(new_n1347), .ZN(G402));
endmodule


