

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  AND2_X1 U322 ( .A1(G229GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U323 ( .A(n368), .B(n367), .ZN(n541) );
  XNOR2_X1 U324 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n359) );
  XNOR2_X1 U325 ( .A(n360), .B(n359), .ZN(n366) );
  XNOR2_X1 U326 ( .A(n333), .B(n290), .ZN(n334) );
  XNOR2_X1 U327 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U328 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n432), .B(n431), .ZN(n450) );
  XOR2_X1 U330 ( .A(n449), .B(n448), .Z(n527) );
  XNOR2_X1 U331 ( .A(n451), .B(KEYINPUT124), .ZN(n452) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(G78GAT), .B(G155GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(G183GAT), .B(G71GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U336 ( .A(n293), .B(G211GAT), .Z(n295) );
  XOR2_X1 U337 ( .A(G15GAT), .B(G1GAT), .Z(n333) );
  XNOR2_X1 U338 ( .A(n333), .B(G127GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n300) );
  XNOR2_X1 U340 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n296), .B(KEYINPUT69), .ZN(n345) );
  XOR2_X1 U342 ( .A(n345), .B(KEYINPUT76), .Z(n298) );
  NAND2_X1 U343 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U346 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n302) );
  XNOR2_X1 U347 ( .A(G22GAT), .B(KEYINPUT15), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n304) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(G64GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U353 ( .A(n308), .B(n307), .Z(n464) );
  XOR2_X1 U354 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n310) );
  XNOR2_X1 U355 ( .A(KEYINPUT75), .B(KEYINPUT66), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(n311), .B(G106GAT), .Z(n313) );
  XOR2_X1 U358 ( .A(G218GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(n413), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .ZN(n314) );
  XOR2_X1 U362 ( .A(n314), .B(G92GAT), .Z(n339) );
  XOR2_X1 U363 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U364 ( .A(n339), .B(n436), .ZN(n316) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U367 ( .A(n318), .B(n317), .Z(n327) );
  INV_X1 U368 ( .A(KEYINPUT7), .ZN(n322) );
  XOR2_X1 U369 ( .A(KEYINPUT8), .B(G50GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G29GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n329) );
  XOR2_X1 U373 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n324) );
  XNOR2_X1 U374 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n329), .B(n325), .ZN(n326) );
  XOR2_X1 U377 ( .A(n327), .B(n326), .Z(n566) );
  INV_X1 U378 ( .A(n566), .ZN(n553) );
  INV_X1 U379 ( .A(n464), .ZN(n582) );
  XOR2_X1 U380 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n328), .B(G8GAT), .ZN(n381) );
  XOR2_X1 U383 ( .A(KEYINPUT30), .B(n381), .Z(n331) );
  XNOR2_X1 U384 ( .A(n329), .B(KEYINPUT29), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n419), .B(n332), .Z(n335) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(G197GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n362) );
  XNOR2_X1 U389 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n353) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n338), .B(G148GAT), .ZN(n412) );
  XNOR2_X1 U392 ( .A(n412), .B(n339), .ZN(n352) );
  XOR2_X1 U393 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n341) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U396 ( .A(n342), .B(KEYINPUT31), .Z(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT70), .B(G64GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n376) );
  XNOR2_X1 U400 ( .A(n345), .B(n376), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U402 ( .A(n348), .B(KEYINPUT71), .Z(n350) );
  XOR2_X1 U403 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U404 ( .A(n435), .B(KEYINPUT72), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n578) );
  XNOR2_X1 U407 ( .A(n353), .B(n578), .ZN(n548) );
  NAND2_X1 U408 ( .A1(n362), .A2(n548), .ZN(n355) );
  INV_X1 U409 ( .A(KEYINPUT46), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  NOR2_X1 U411 ( .A1(n582), .A2(n356), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n357), .B(KEYINPUT115), .ZN(n358) );
  NOR2_X1 U413 ( .A1(n553), .A2(n358), .ZN(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT36), .B(n566), .Z(n584) );
  NAND2_X1 U415 ( .A1(n582), .A2(n584), .ZN(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT45), .B(n361), .Z(n364) );
  XNOR2_X1 U417 ( .A(KEYINPUT68), .B(n362), .ZN(n530) );
  NOR2_X1 U418 ( .A1(n530), .A2(n578), .ZN(n363) );
  NAND2_X1 U419 ( .A1(n364), .A2(n363), .ZN(n365) );
  NAND2_X1 U420 ( .A1(n366), .A2(n365), .ZN(n368) );
  XNOR2_X1 U421 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n367) );
  XOR2_X1 U422 ( .A(G92GAT), .B(G218GAT), .Z(n370) );
  NAND2_X1 U423 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(KEYINPUT96), .B(n371), .Z(n375) );
  XOR2_X1 U426 ( .A(G183GAT), .B(KEYINPUT17), .Z(n373) );
  XNOR2_X1 U427 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n440) );
  XNOR2_X1 U429 ( .A(n440), .B(G190GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U431 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(n380), .ZN(n428) );
  XOR2_X1 U436 ( .A(n381), .B(n428), .Z(n382) );
  XOR2_X1 U437 ( .A(n383), .B(n382), .Z(n500) );
  INV_X1 U438 ( .A(n500), .ZN(n518) );
  NAND2_X1 U439 ( .A1(n541), .A2(n518), .ZN(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n573) );
  XOR2_X1 U442 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n387) );
  XNOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U445 ( .A(KEYINPUT95), .B(G57GAT), .Z(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n403) );
  XOR2_X1 U449 ( .A(KEYINPUT0), .B(G127GAT), .Z(n393) );
  XNOR2_X1 U450 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U452 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n394) );
  XOR2_X1 U453 ( .A(n395), .B(n394), .Z(n449) );
  INV_X1 U454 ( .A(n449), .ZN(n401) );
  XOR2_X1 U455 ( .A(G155GAT), .B(KEYINPUT88), .Z(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n423) );
  XOR2_X1 U458 ( .A(n423), .B(KEYINPUT94), .Z(n399) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U461 ( .A(n401), .B(n400), .Z(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n411) );
  XOR2_X1 U463 ( .A(KEYINPUT91), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(G1GAT), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U466 ( .A(G162GAT), .B(G120GAT), .Z(n407) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G134GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U469 ( .A(n409), .B(n408), .Z(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n513) );
  XNOR2_X1 U471 ( .A(G85GAT), .B(n513), .ZN(n468) );
  INV_X1 U472 ( .A(n468), .ZN(n572) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U476 ( .A(G204GAT), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT90), .B(KEYINPUT85), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(n418), .B(KEYINPUT22), .Z(n421) );
  XNOR2_X1 U480 ( .A(G50GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U482 ( .A(n422), .B(KEYINPUT89), .Z(n425) );
  XNOR2_X1 U483 ( .A(n423), .B(KEYINPUT24), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n461) );
  AND2_X1 U487 ( .A1(n572), .A2(n461), .ZN(n430) );
  NAND2_X1 U488 ( .A1(n573), .A2(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(KEYINPUT20), .B(G176GAT), .Z(n434) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U492 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n438) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n439), .B(G99GAT), .Z(n445) );
  XOR2_X1 U496 ( .A(G15GAT), .B(n440), .Z(n442) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n448) );
  NAND2_X1 U502 ( .A1(n450), .A2(n527), .ZN(n565) );
  NOR2_X1 U503 ( .A1(n464), .A2(n565), .ZN(n453) );
  INV_X1 U504 ( .A(G183GAT), .ZN(n451) );
  INV_X1 U505 ( .A(n530), .ZN(n556) );
  NOR2_X1 U506 ( .A1(n556), .A2(n578), .ZN(n483) );
  NAND2_X1 U507 ( .A1(n527), .A2(n518), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n461), .A2(n454), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT25), .ZN(n458) );
  NOR2_X1 U510 ( .A1(n461), .A2(n527), .ZN(n456) );
  XOR2_X1 U511 ( .A(n456), .B(KEYINPUT26), .Z(n542) );
  XNOR2_X1 U512 ( .A(n500), .B(KEYINPUT27), .ZN(n460) );
  NOR2_X1 U513 ( .A1(n542), .A2(n460), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n458), .A2(n457), .ZN(n459) );
  NOR2_X1 U515 ( .A1(n468), .A2(n459), .ZN(n463) );
  NOR2_X1 U516 ( .A1(n460), .A2(n572), .ZN(n543) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n461), .Z(n522) );
  INV_X1 U518 ( .A(n522), .ZN(n507) );
  NAND2_X1 U519 ( .A1(n543), .A2(n507), .ZN(n529) );
  NOR2_X1 U520 ( .A1(n527), .A2(n529), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n480) );
  NOR2_X1 U522 ( .A1(n553), .A2(n464), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n465), .Z(n466) );
  NOR2_X1 U524 ( .A1(n480), .A2(n466), .ZN(n496) );
  NAND2_X1 U525 ( .A1(n483), .A2(n496), .ZN(n467) );
  XNOR2_X1 U526 ( .A(KEYINPUT97), .B(n467), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n476), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(KEYINPUT34), .ZN(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  NAND2_X1 U530 ( .A1(n476), .A2(n518), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U532 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n473) );
  NAND2_X1 U533 ( .A1(n476), .A2(n527), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(n475) );
  XOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT98), .Z(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n478) );
  NAND2_X1 U538 ( .A1(n476), .A2(n522), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(n479), .ZN(G1327GAT) );
  NOR2_X1 U541 ( .A1(n582), .A2(n480), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n481), .A2(n584), .ZN(n482) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n482), .ZN(n512) );
  NAND2_X1 U544 ( .A1(n483), .A2(n512), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT38), .ZN(n493) );
  NOR2_X1 U546 ( .A1(n493), .A2(n572), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n493), .A2(n500), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1329GAT) );
  INV_X1 U553 ( .A(n527), .ZN(n503) );
  NOR2_X1 U554 ( .A1(n493), .A2(n503), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n492), .Z(G1330GAT) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n495) );
  NOR2_X1 U559 ( .A1(n507), .A2(n493), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  XNOR2_X1 U561 ( .A(KEYINPUT107), .B(n548), .ZN(n560) );
  NOR2_X1 U562 ( .A1(n362), .A2(n560), .ZN(n511) );
  NAND2_X1 U563 ( .A1(n511), .A2(n496), .ZN(n506) );
  NOR2_X1 U564 ( .A1(n572), .A2(n506), .ZN(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U566 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n499), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n500), .A2(n506), .ZN(n501) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n501), .Z(n502) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n503), .A2(n506), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  AND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n523) );
  OR2_X1 U579 ( .A1(G85GAT), .A2(n523), .ZN(n515) );
  NAND2_X1 U580 ( .A1(n523), .A2(n513), .ZN(n514) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT111), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT113), .Z(n520) );
  NAND2_X1 U585 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n527), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n541), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n538), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  INV_X1 U597 ( .A(n538), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n560), .A2(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U602 ( .A1(n538), .A2(n582), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n553), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n547) );
  INV_X1 U609 ( .A(n541), .ZN(n545) );
  INV_X1 U610 ( .A(n542), .ZN(n574) );
  NAND2_X1 U611 ( .A1(n543), .A2(n574), .ZN(n544) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n362), .A2(n554), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n582), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n565), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT122), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n565), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  INV_X1 U633 ( .A(G190GAT), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT58), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n577) );
  AND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  AND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n362), .ZN(n576) );
  XOR2_X1 U642 ( .A(n577), .B(n576), .Z(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

