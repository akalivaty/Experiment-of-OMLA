//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT28), .Z(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT68), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n211), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n223), .B2(new_n220), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n216), .A2(new_n218), .A3(new_n219), .A4(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n214), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n229), .A2(KEYINPUT69), .B1(G127gat), .B2(G134gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G127gat), .B2(G134gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n228), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n211), .A2(new_n235), .A3(KEYINPUT67), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(new_n236), .C1(G183gat), .C2(G190gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n211), .B(KEYINPUT66), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n206), .A3(new_n217), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT25), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n214), .A3(new_n225), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT33), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(KEYINPUT32), .ZN(new_n251));
  XOR2_X1   g050(.A(G15gat), .B(G43gat), .Z(new_n252));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT34), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n254), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n248), .B(KEYINPUT32), .C1(new_n249), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n255), .A2(new_n258), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n258), .B1(new_n255), .B2(new_n260), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT36), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT36), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n262), .B2(new_n264), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(KEYINPUT71), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  INV_X1    g075(.A(G218gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(KEYINPUT22), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT72), .ZN(new_n280));
  XOR2_X1   g079(.A(G211gat), .B(G218gat), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n283), .A3(KEYINPUT72), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT73), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n243), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n226), .B2(new_n241), .ZN(new_n289));
  INV_X1    g088(.A(new_n286), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n285), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n285), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n243), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n286), .B1(new_n226), .B2(new_n241), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n291), .A2(new_n296), .A3(KEYINPUT30), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n291), .A2(new_n296), .A3(new_n300), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n296), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n299), .B(KEYINPUT74), .Z(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G1gat), .B(G29gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(KEYINPUT77), .B1(KEYINPUT2), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(KEYINPUT77), .B2(new_n323), .ZN(new_n326));
  XOR2_X1   g125(.A(G155gat), .B(G162gat), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT79), .B(G155gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G162gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT78), .B(G141gat), .Z(new_n333));
  OAI21_X1  g132(.A(new_n322), .B1(new_n333), .B2(new_n320), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n328), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n232), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n331), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT80), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n343), .A2(new_n335), .B1(new_n327), .B2(new_n326), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n233), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n232), .B(KEYINPUT81), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n328), .B(new_n350), .C1(new_n336), .C2(new_n337), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(G225gat), .A3(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT39), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n338), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n356), .A2(new_n345), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n319), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(KEYINPUT39), .B2(new_n354), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT40), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n356), .B2(new_n345), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(KEYINPUT83), .B(KEYINPUT5), .C1(new_n357), .C2(new_n358), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n341), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n358), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n367), .B(new_n368), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n347), .A2(new_n366), .A3(new_n352), .A4(new_n358), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n361), .A2(new_n362), .B1(new_n376), .B2(new_n319), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n313), .A2(new_n363), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n319), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n318), .A3(new_n375), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n319), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n285), .B1(new_n294), .B2(new_n295), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(KEYINPUT37), .C1(new_n385), .C2(new_n285), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT37), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n291), .A2(new_n296), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT38), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .A4(new_n310), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n306), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n300), .B1(new_n309), .B2(KEYINPUT37), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n389), .B1(new_n392), .B2(new_n388), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n383), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n378), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n285), .B1(new_n351), .B2(new_n293), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n279), .B(new_n281), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n400), .B2(new_n293), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n344), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n282), .A2(new_n293), .A3(new_n284), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n350), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n398), .B1(new_n338), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n344), .B2(new_n350), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(new_n285), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n403), .B2(new_n408), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n397), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n418), .A2(KEYINPUT87), .A3(new_n413), .A4(new_n410), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n410), .A2(KEYINPUT85), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n408), .A3(new_n422), .A4(new_n409), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(new_n418), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425));
  INV_X1    g224(.A(new_n413), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT88), .B(new_n420), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n274), .B1(new_n396), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT89), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n382), .A2(new_n383), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n435), .B(new_n437), .C1(new_n438), .C2(new_n313), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n313), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n272), .A2(new_n442), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT90), .B(new_n266), .C1(new_n262), .C2(new_n264), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n446));
  NAND4_X1  g245(.A1(new_n441), .A2(new_n445), .A3(new_n433), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n382), .A2(new_n383), .ZN(new_n448));
  INV_X1    g247(.A(new_n313), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n448), .A3(new_n449), .A4(new_n272), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n440), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT101), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OR2_X1    g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458));
  AND2_X1   g257(.A1(G71gat), .A2(G78gat), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(KEYINPUT9), .ZN(new_n460));
  XOR2_X1   g259(.A(G71gat), .B(G78gat), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT100), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(KEYINPUT100), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(G231gat), .A3(G233gat), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G231gat), .A2(G233gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n467), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G127gat), .B(G155gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n472), .A2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n456), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n475), .A3(new_n455), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(G1gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n484));
  AOI21_X1  g283(.A(G8gat), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n485), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n462), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(KEYINPUT21), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n492), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n480), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G183gat), .B(G211gat), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT13), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR3_X1    g309(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(KEYINPUT94), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n515), .B1(new_n510), .B2(new_n511), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n520), .C1(KEYINPUT94), .C2(new_n522), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n490), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n489), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n505), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT96), .B1(new_n529), .B2(KEYINPUT17), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n535), .B(new_n532), .C1(new_n524), .C2(new_n526), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n489), .B(new_n533), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n503), .A3(new_n528), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT11), .ZN(new_n542));
  INV_X1    g341(.A(G169gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT12), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n503), .A4(new_n528), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(KEYINPUT97), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(KEYINPUT97), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n540), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n540), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  INV_X1    g351(.A(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(KEYINPUT98), .A3(new_n553), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT102), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(G99gat), .B2(G106gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(KEYINPUT102), .C1(new_n568), .C2(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT103), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n568), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n568), .A2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n575), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n570), .B2(new_n577), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n582), .B(new_n533), .C1(new_n534), .C2(new_n536), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  AND2_X1   g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n527), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n588), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n583), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n589), .B2(new_n593), .ZN(new_n595));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596));
  OR3_X1    g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n596), .B1(new_n594), .B2(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n491), .B1(new_n580), .B2(new_n581), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n570), .A2(new_n577), .ZN(new_n603));
  INV_X1    g402(.A(new_n579), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n462), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(KEYINPUT10), .B(new_n491), .C1(new_n580), .C2(new_n581), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT104), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT104), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n601), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n600), .B1(new_n602), .B2(new_n607), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n619), .B(KEYINPUT105), .Z(new_n622));
  AOI21_X1  g421(.A(new_n601), .B1(new_n609), .B2(new_n610), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(new_n616), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n624), .A2(KEYINPUT106), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(KEYINPUT106), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR4_X1   g426(.A1(new_n502), .A2(new_n558), .A3(new_n599), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n453), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n448), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n449), .ZN(new_n632));
  INV_X1    g431(.A(G8gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT42), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT16), .B(G8gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  MUX2_X1   g435(.A(KEYINPUT42), .B(new_n634), .S(new_n636), .Z(G1325gat));
  INV_X1    g436(.A(new_n274), .ZN(new_n638));
  OAI21_X1  g437(.A(G15gat), .B1(new_n629), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n445), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(G15gat), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n629), .B2(new_n641), .ZN(G1326gat));
  NAND2_X1  g441(.A1(new_n435), .A2(new_n437), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  AND2_X1   g445(.A1(new_n597), .A2(new_n598), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n440), .B2(new_n452), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n501), .A2(new_n558), .A3(new_n627), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G29gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n438), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT45), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n434), .A2(new_n439), .B1(new_n447), .B2(new_n451), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n647), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n649), .ZN(new_n659));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659), .B2(new_n448), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n660), .ZN(G1328gat));
  INV_X1    g460(.A(G36gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n650), .A2(new_n662), .A3(new_n313), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT46), .Z(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n659), .B2(new_n449), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n654), .A2(new_n657), .A3(new_n274), .A4(new_n649), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G43gat), .ZN(new_n669));
  INV_X1    g468(.A(G43gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n650), .A2(new_n670), .A3(new_n445), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1330gat));
  INV_X1    g473(.A(G50gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n659), .ZN(new_n676));
  INV_X1    g475(.A(new_n433), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n643), .A2(G50gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n650), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT48), .ZN(new_n681));
  INV_X1    g480(.A(new_n643), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n658), .A2(new_n682), .A3(new_n649), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n683), .A2(G50gat), .B1(new_n650), .B2(new_n679), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n678), .A2(new_n681), .B1(new_n684), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g484(.A(new_n627), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n501), .A2(new_n558), .A3(new_n647), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n656), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n438), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g489(.A(new_n449), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT108), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1333gat));
  NAND3_X1  g494(.A1(new_n688), .A2(G71gat), .A3(new_n274), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n688), .A2(new_n445), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G71gat), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n688), .A2(new_n682), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  AND3_X1   g501(.A1(new_n552), .A2(KEYINPUT98), .A3(new_n553), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT98), .B1(new_n552), .B2(new_n553), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n550), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n501), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n648), .A2(KEYINPUT51), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT51), .B1(new_n648), .B2(new_n706), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n709), .A2(new_n564), .A3(new_n438), .A4(new_n627), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n654), .A2(new_n657), .A3(new_n627), .A4(new_n706), .ZN(new_n711));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711), .B2(new_n448), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1336gat));
  AND3_X1   g512(.A1(new_n654), .A2(new_n657), .A3(new_n706), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n313), .A4(new_n627), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT110), .B1(new_n711), .B2(new_n449), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n565), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n449), .A2(new_n686), .A3(G92gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n707), .B2(new_n708), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G92gat), .B1(new_n711), .B2(new_n449), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(new_n720), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n718), .A2(new_n722), .B1(new_n724), .B2(new_n721), .ZN(G1337gat));
  NOR3_X1   g524(.A1(new_n640), .A2(G99gat), .A3(new_n686), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G99gat), .B1(new_n711), .B2(new_n638), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1338gat));
  NOR3_X1   g528(.A1(new_n433), .A2(G106gat), .A3(new_n686), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n707), .B2(new_n708), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n732));
  OAI21_X1  g531(.A(G106gat), .B1(new_n711), .B2(new_n643), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n730), .C1(new_n707), .C2(new_n708), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT53), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT53), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n433), .A2(new_n686), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n654), .A2(new_n657), .A3(new_n706), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT112), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G106gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(KEYINPUT112), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n738), .B(new_n731), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(G1339gat));
  AND4_X1   g544(.A1(new_n558), .A2(new_n501), .A3(new_n647), .A4(new_n686), .ZN(new_n746));
  INV_X1    g545(.A(new_n619), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n623), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n609), .A2(new_n610), .A3(new_n601), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT54), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n615), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT55), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(new_n749), .C1(new_n615), .C2(new_n751), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n620), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n528), .A2(new_n530), .A3(new_n505), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT113), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n528), .A2(new_n759), .A3(new_n530), .A4(new_n505), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n503), .B1(new_n537), .B2(new_n528), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n545), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n765), .B(new_n545), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n599), .A2(new_n550), .A3(new_n756), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(new_n627), .A3(new_n550), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n705), .B2(new_n756), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n771), .B2(new_n599), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n746), .B1(new_n772), .B2(new_n502), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n682), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n438), .A2(new_n449), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n640), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(G113gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n558), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n773), .A2(new_n448), .A3(new_n677), .A4(new_n268), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n449), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n705), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n778), .ZN(G1340gat));
  INV_X1    g582(.A(G120gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n777), .A2(new_n784), .A3(new_n686), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n627), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n784), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT115), .Z(G1341gat));
  INV_X1    g587(.A(G127gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n781), .A2(new_n789), .A3(new_n501), .ZN(new_n790));
  OAI21_X1  g589(.A(G127gat), .B1(new_n777), .B2(new_n502), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1342gat));
  NAND2_X1  g591(.A1(new_n449), .A2(new_n599), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(G134gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT56), .Z(new_n796));
  OAI21_X1  g595(.A(G134gat), .B1(new_n777), .B2(new_n647), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1343gat));
  NOR2_X1   g601(.A1(new_n274), .A2(new_n775), .ZN(new_n803));
  INV_X1    g602(.A(new_n746), .ZN(new_n804));
  INV_X1    g603(.A(new_n768), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n753), .A2(new_n755), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n806), .B2(new_n621), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n808), .B(new_n620), .C1(new_n753), .C2(new_n755), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n769), .B1(new_n558), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n805), .B1(new_n811), .B2(new_n647), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n812), .B2(new_n501), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT57), .A4(new_n682), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n773), .B2(new_n433), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n755), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n613), .B1(new_n609), .B2(new_n610), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n600), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n751), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n754), .B1(new_n824), .B2(new_n749), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n621), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n808), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n756), .A2(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n770), .B1(new_n705), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n768), .B1(new_n830), .B2(new_n599), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n502), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n643), .B1(new_n832), .B2(new_n804), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n814), .B1(new_n833), .B2(KEYINPUT57), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n705), .B(new_n803), .C1(new_n818), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n333), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT119), .B1(new_n773), .B2(new_n448), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n769), .B1(new_n558), .B2(new_n826), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n647), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n501), .B1(new_n840), .B2(new_n768), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n838), .B(new_n438), .C1(new_n841), .C2(new_n746), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n274), .A2(new_n433), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n449), .A2(new_n837), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n558), .A2(G141gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n836), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT58), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n836), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(KEYINPUT120), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  AOI221_X4 g651(.A(KEYINPUT58), .B1(new_n844), .B2(new_n845), .C1(new_n835), .C2(new_n333), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n849), .B1(new_n836), .B2(new_n846), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(G1344gat));
  NAND3_X1  g655(.A1(new_n844), .A2(new_n320), .A3(new_n627), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT121), .Z(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n803), .B(KEYINPUT122), .Z(new_n860));
  OR2_X1    g659(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n677), .C1(new_n841), .C2(new_n746), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n686), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n320), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n627), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT123), .B1(new_n867), .B2(new_n860), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n859), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n803), .B1(new_n818), .B2(new_n834), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(new_n686), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n871), .A2(new_n859), .A3(G148gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n858), .B1(new_n869), .B2(new_n872), .ZN(G1345gat));
  OAI21_X1  g672(.A(new_n329), .B1(new_n870), .B2(new_n502), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n502), .A2(new_n329), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n844), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n870), .B2(new_n647), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n793), .A2(G162gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n837), .A2(new_n842), .A3(new_n843), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n438), .A2(new_n449), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n774), .A2(new_n445), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(G169gat), .A3(new_n705), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n773), .A2(new_n438), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n677), .A2(new_n449), .A3(new_n268), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n543), .B1(new_n887), .B2(new_n558), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(G1348gat));
  NAND3_X1  g689(.A1(new_n883), .A2(G176gat), .A3(new_n627), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n887), .A2(new_n686), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(G176gat), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT125), .Z(G1349gat));
  NAND2_X1  g693(.A1(new_n883), .A2(new_n501), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G183gat), .ZN(new_n896));
  INV_X1    g695(.A(new_n887), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n501), .A2(new_n202), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n897), .A2(new_n898), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n900), .B(new_n901), .Z(G1350gat));
  AOI21_X1  g701(.A(new_n203), .B1(new_n883), .B2(new_n599), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT61), .Z(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n203), .A3(new_n599), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1351gat));
  NAND2_X1  g705(.A1(new_n843), .A2(new_n313), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT127), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n885), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n705), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n638), .A2(new_n882), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n861), .B2(new_n862), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n705), .A2(G197gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  NOR3_X1   g714(.A1(new_n909), .A2(G204gat), .A3(new_n686), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT62), .ZN(new_n917));
  OAI21_X1  g716(.A(G204gat), .B1(new_n867), .B2(new_n912), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n910), .A2(new_n276), .A3(new_n501), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n913), .A2(new_n501), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  NAND3_X1  g723(.A1(new_n910), .A2(new_n277), .A3(new_n599), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n913), .A2(new_n599), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n277), .ZN(G1355gat));
endmodule


