

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U326 ( .A(n418), .B(KEYINPUT64), .ZN(n573) );
  INV_X1 U327 ( .A(KEYINPUT15), .ZN(n305) );
  XNOR2_X1 U328 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U329 ( .A(KEYINPUT41), .B(n578), .Z(n557) );
  AND2_X1 U330 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U331 ( .A(n383), .B(n321), .Z(n295) );
  AND2_X1 U332 ( .A1(n574), .A2(n557), .ZN(n344) );
  NOR2_X1 U333 ( .A1(n533), .A2(n392), .ZN(n393) );
  XNOR2_X1 U334 ( .A(n334), .B(n294), .ZN(n335) );
  XNOR2_X1 U335 ( .A(n336), .B(n335), .ZN(n341) );
  XNOR2_X1 U336 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U337 ( .A(n314), .B(n313), .Z(n544) );
  XNOR2_X1 U338 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U339 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT12), .B(KEYINPUT82), .Z(n297) );
  XNOR2_X1 U341 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n314) );
  XOR2_X1 U343 ( .A(G64GAT), .B(KEYINPUT14), .Z(n299) );
  XNOR2_X1 U344 ( .A(G1GAT), .B(G57GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U346 ( .A(G78GAT), .B(G211GAT), .Z(n301) );
  XNOR2_X1 U347 ( .A(G127GAT), .B(G155GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n312) );
  XNOR2_X1 U350 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n304) );
  XOR2_X1 U351 ( .A(n304), .B(KEYINPUT13), .Z(n331) );
  XOR2_X1 U352 ( .A(n331), .B(KEYINPUT79), .Z(n306) );
  XOR2_X1 U353 ( .A(G8GAT), .B(G183GAT), .Z(n383) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G22GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(KEYINPUT69), .ZN(n321) );
  NAND2_X1 U356 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n295), .B(n308), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  INV_X1 U359 ( .A(n544), .ZN(n582) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G36GAT), .Z(n316) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G50GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U363 ( .A(KEYINPUT68), .B(G8GAT), .Z(n318) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(G197GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n329) );
  XOR2_X1 U367 ( .A(G113GAT), .B(G1GAT), .Z(n412) );
  XOR2_X1 U368 ( .A(n412), .B(n321), .Z(n323) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(n324), .B(KEYINPUT30), .Z(n327) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n325), .B(KEYINPUT7), .ZN(n360) );
  XNOR2_X1 U374 ( .A(n360), .B(KEYINPUT29), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U376 ( .A(n329), .B(n328), .Z(n574) );
  XNOR2_X1 U377 ( .A(G99GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n330), .B(KEYINPUT73), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n349), .B(n331), .ZN(n343) );
  XOR2_X1 U380 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G57GAT), .Z(n408) );
  XOR2_X1 U382 ( .A(n387), .B(n408), .Z(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n333) );
  XNOR2_X1 U384 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U386 ( .A(KEYINPUT72), .B(G78GAT), .Z(n421) );
  XOR2_X1 U387 ( .A(G92GAT), .B(G85GAT), .Z(n338) );
  XNOR2_X1 U388 ( .A(G148GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n421), .B(n339), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n578) );
  XNOR2_X1 U393 ( .A(n344), .B(KEYINPUT46), .ZN(n345) );
  NOR2_X1 U394 ( .A1(n582), .A2(n345), .ZN(n346) );
  XNOR2_X1 U395 ( .A(n346), .B(KEYINPUT114), .ZN(n365) );
  XOR2_X1 U396 ( .A(G92GAT), .B(G218GAT), .Z(n348) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(G190GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n380) );
  XNOR2_X1 U399 ( .A(n380), .B(n349), .ZN(n364) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  XOR2_X1 U401 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n351) );
  XNOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT67), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U404 ( .A(n420), .B(n352), .Z(n354) );
  NAND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n356) );
  XNOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT9), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n362) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G134GAT), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n359), .B(G85GAT), .ZN(n398) );
  XOR2_X1 U413 ( .A(n360), .B(n398), .Z(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n563) );
  NAND2_X1 U416 ( .A1(n365), .A2(n563), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n366), .B(KEYINPUT115), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n367), .B(KEYINPUT47), .ZN(n375) );
  XNOR2_X1 U419 ( .A(KEYINPUT116), .B(KEYINPUT45), .ZN(n370) );
  INV_X1 U420 ( .A(KEYINPUT78), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n563), .B(n368), .ZN(n458) );
  XOR2_X1 U422 ( .A(KEYINPUT36), .B(n458), .Z(n587) );
  NOR2_X1 U423 ( .A1(n544), .A2(n587), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(n371), .B(KEYINPUT66), .Z(n372) );
  NOR2_X1 U426 ( .A1(n578), .A2(n372), .ZN(n373) );
  INV_X1 U427 ( .A(n574), .ZN(n538) );
  NAND2_X1 U428 ( .A1(n373), .A2(n538), .ZN(n374) );
  NAND2_X1 U429 ( .A1(n374), .A2(n375), .ZN(n377) );
  XNOR2_X1 U430 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n533) );
  XOR2_X1 U432 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n379) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n438) );
  XNOR2_X1 U435 ( .A(n438), .B(n380), .ZN(n391) );
  XOR2_X1 U436 ( .A(G204GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n419) );
  XOR2_X1 U439 ( .A(n383), .B(n419), .Z(n385) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(n386), .B(KEYINPUT95), .Z(n389) );
  XNOR2_X1 U443 ( .A(n387), .B(KEYINPUT96), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(n391), .B(n390), .Z(n495) );
  XOR2_X1 U446 ( .A(n495), .B(KEYINPUT123), .Z(n392) );
  XNOR2_X1 U447 ( .A(KEYINPUT54), .B(n393), .ZN(n417) );
  XNOR2_X1 U448 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(KEYINPUT2), .ZN(n395) );
  XOR2_X1 U450 ( .A(n395), .B(KEYINPUT87), .Z(n397) );
  XNOR2_X1 U451 ( .A(G141GAT), .B(G148GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n433) );
  XOR2_X1 U453 ( .A(n398), .B(KEYINPUT92), .Z(n400) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n433), .B(n401), .ZN(n416) );
  XOR2_X1 U457 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT88), .B(KEYINPUT93), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U460 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n405) );
  XNOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT90), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n407), .B(n406), .Z(n414) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(n408), .Z(n410) );
  XOR2_X1 U465 ( .A(KEYINPUT0), .B(G127GAT), .Z(n437) );
  XNOR2_X1 U466 ( .A(n437), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n472) );
  XOR2_X1 U471 ( .A(KEYINPUT94), .B(n472), .Z(n520) );
  INV_X1 U472 ( .A(n520), .ZN(n490) );
  NAND2_X1 U473 ( .A1(n417), .A2(n490), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n424) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n431) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(G106GAT), .Z(n428) );
  XNOR2_X1 U481 ( .A(G22GAT), .B(G218GAT), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n429), .B(KEYINPUT24), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n466) );
  NOR2_X1 U486 ( .A1(n573), .A2(n466), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n434), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U488 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G134GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n440) );
  XNOR2_X1 U492 ( .A(G190GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U494 ( .A(G71GAT), .B(G183GAT), .Z(n442) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U498 ( .A(G120GAT), .B(G176GAT), .Z(n446) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(KEYINPUT85), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(G113GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U503 ( .A(n451), .B(n450), .Z(n534) );
  INV_X1 U504 ( .A(n534), .ZN(n499) );
  NOR2_X2 U505 ( .A1(n452), .A2(n499), .ZN(n567) );
  NAND2_X1 U506 ( .A1(n567), .A2(n557), .ZN(n456) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U508 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n578), .A2(n538), .ZN(n457) );
  XOR2_X1 U510 ( .A(n457), .B(KEYINPUT74), .Z(n488) );
  INV_X1 U511 ( .A(n458), .ZN(n548) );
  NAND2_X1 U512 ( .A1(n548), .A2(n582), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT83), .ZN(n475) );
  XNOR2_X1 U515 ( .A(KEYINPUT28), .B(n466), .ZN(n527) );
  XOR2_X1 U516 ( .A(n495), .B(KEYINPUT27), .Z(n468) );
  NAND2_X1 U517 ( .A1(n520), .A2(n468), .ZN(n532) );
  NOR2_X1 U518 ( .A1(n527), .A2(n532), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT97), .B(n461), .Z(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n499), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT98), .ZN(n474) );
  NOR2_X1 U522 ( .A1(n499), .A2(n495), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n466), .A2(n464), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT25), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n466), .A2(n499), .ZN(n467) );
  XOR2_X1 U526 ( .A(n467), .B(KEYINPUT26), .Z(n571) );
  NAND2_X1 U527 ( .A1(n468), .A2(n571), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n485) );
  NAND2_X1 U531 ( .A1(n475), .A2(n485), .ZN(n505) );
  NOR2_X1 U532 ( .A1(n488), .A2(n505), .ZN(n481) );
  NAND2_X1 U533 ( .A1(n520), .A2(n481), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  INV_X1 U536 ( .A(n495), .ZN(n522) );
  NAND2_X1 U537 ( .A1(n481), .A2(n522), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n534), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n483) );
  NAND2_X1 U543 ( .A1(n481), .A2(n527), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n544), .A2(n485), .ZN(n486) );
  NOR2_X1 U547 ( .A1(n587), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n487), .ZN(n519) );
  OR2_X1 U549 ( .A1(n488), .A2(n519), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT38), .ZN(n503) );
  NOR2_X1 U551 ( .A1(n490), .A2(n503), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n503), .A2(n495), .ZN(n497) );
  XNOR2_X1 U557 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NOR2_X1 U560 ( .A1(n503), .A2(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  INV_X1 U564 ( .A(n527), .ZN(n536) );
  NOR2_X1 U565 ( .A1(n503), .A2(n536), .ZN(n504) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n508) );
  NAND2_X1 U568 ( .A1(n557), .A2(n538), .ZN(n518) );
  NOR2_X1 U569 ( .A1(n518), .A2(n505), .ZN(n506) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(n506), .Z(n513) );
  NAND2_X1 U571 ( .A1(n513), .A2(n520), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n522), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT108), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n534), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U580 ( .A1(n513), .A2(n527), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT110), .Z(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n520), .A2(n528), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT111), .Z(n524) );
  NAND2_X1 U588 ( .A1(n528), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n534), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT112), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n530) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n551) );
  NAND2_X1 U598 ( .A1(n534), .A2(n551), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(n535), .Z(n537) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n538), .A2(n547), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(KEYINPUT119), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  INV_X1 U604 ( .A(n557), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n541), .A2(n547), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n544), .A2(n547), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n571), .A2(n551), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT120), .B(n552), .ZN(n562) );
  INV_X1 U616 ( .A(n562), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n574), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(n556), .Z(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n582), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n567), .A2(n574), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n582), .A2(n567), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n458), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  INV_X1 U638 ( .A(n571), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U640 ( .A1(n585), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(KEYINPUT62), .ZN(n589) );
  INV_X1 U651 ( .A(n585), .ZN(n586) );
  NOR2_X1 U652 ( .A1(n586), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

