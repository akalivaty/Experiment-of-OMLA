//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G97), .A2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G58), .C2(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n228), .A2(new_n217), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  INV_X1    g0036(.A(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n208), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n207), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n254), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n217), .A2(new_n253), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n259), .B1(new_n258), .B2(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n229), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n202), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n264), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n216), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G50), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT9), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n280), .B1(new_n281), .B2(new_n278), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT67), .B1(new_n253), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n229), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G33), .A3(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n275), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n286), .B1(new_n237), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n274), .A2(new_n296), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n272), .C1(G179), .C2(new_n294), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(G58), .B(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(G159), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n261), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT3), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT7), .B(new_n217), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(G20), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT77), .B1(new_n320), .B2(KEYINPUT7), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT7), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT77), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(new_n278), .C2(G20), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n317), .A2(new_n321), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n327), .A2(KEYINPUT79), .A3(G68), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT79), .B1(new_n327), .B2(G68), .ZN(new_n329));
  OAI211_X1 g0129(.A(KEYINPUT16), .B(new_n312), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT80), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n313), .B2(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n253), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n319), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n325), .B1(new_n278), .B2(G20), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n212), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n331), .B1(new_n338), .B2(new_n311), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n264), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n278), .A2(G223), .A3(new_n279), .ZN(new_n341));
  INV_X1    g0141(.A(G87), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(new_n253), .B2(new_n342), .C1(new_n282), .C2(new_n237), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n277), .B1(new_n343), .B2(new_n285), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n292), .A2(G232), .A3(new_n275), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  INV_X1    g0147(.A(new_n269), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n256), .A2(new_n270), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(new_n266), .B2(new_n256), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(G190), .A3(new_n345), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n340), .A2(new_n347), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT17), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n344), .A2(G179), .A3(new_n345), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n303), .B1(new_n344), .B2(new_n345), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n340), .B2(new_n351), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT81), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n318), .A2(new_n319), .A3(G226), .A4(new_n279), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n318), .A2(new_n319), .A3(G232), .A4(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n285), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n292), .A2(G238), .A3(new_n275), .ZN(new_n371));
  INV_X1    g0171(.A(new_n277), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n370), .A2(new_n376), .A3(new_n371), .A4(new_n372), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  OR3_X1    g0178(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT13), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(G200), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n374), .A2(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G190), .ZN(new_n382));
  INV_X1    g0182(.A(new_n264), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT70), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(new_n216), .A3(G13), .A4(G20), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n383), .A2(new_n384), .A3(new_n270), .A4(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n212), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT12), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n212), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n212), .A2(G20), .ZN(new_n393));
  OR4_X1    g0193(.A1(KEYINPUT12), .A2(new_n393), .A3(G1), .A4(new_n223), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n254), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n393), .B1(new_n202), .B2(new_n261), .C1(new_n396), .C2(new_n281), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n264), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT11), .Z(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n380), .A2(new_n382), .A3(new_n395), .A4(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n307), .A2(new_n354), .A3(new_n365), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n378), .A2(new_n379), .A3(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n381), .A2(G179), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n378), .A2(new_n379), .A3(G169), .A4(new_n404), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n400), .A2(new_n395), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n406), .A2(KEYINPUT76), .A3(new_n407), .A4(new_n408), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n390), .A2(new_n281), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT71), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n255), .A2(new_n261), .B1(new_n217), .B2(new_n281), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n396), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n264), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT72), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n387), .A2(new_n281), .ZN(new_n423));
  OR3_X1    g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n421), .B2(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G244), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n372), .B1(new_n293), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n278), .A2(G232), .A3(new_n279), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(new_n249), .B2(new_n278), .C1(new_n282), .C2(new_n213), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n285), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n429), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n303), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  INV_X1    g0237(.A(G179), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n426), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(G190), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(G200), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n424), .A3(new_n425), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n414), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n402), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G294), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n318), .A2(new_n319), .A3(G250), .A4(new_n279), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n285), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G264), .A3(new_n292), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n454), .A2(KEYINPUT82), .A3(G274), .A4(new_n456), .ZN(new_n461));
  INV_X1    g0261(.A(new_n453), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n456), .B(G274), .C1(new_n462), .C2(new_n451), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n303), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT90), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n469), .A3(new_n458), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n450), .B2(new_n458), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n473), .B2(new_n438), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n318), .A2(new_n319), .A3(new_n217), .A4(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT88), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT88), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n278), .A2(new_n477), .A3(new_n217), .A4(G87), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT22), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n217), .A2(G107), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT23), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT22), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(KEYINPUT88), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n254), .A2(G116), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n479), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(new_n484), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n481), .A4(new_n479), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n383), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n216), .A2(G33), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n269), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n249), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n266), .A2(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT89), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT25), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n474), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n249), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n249), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n217), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n336), .A2(new_n337), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n261), .A2(new_n281), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n264), .B1(new_n500), .B2(new_n267), .ZN(new_n511));
  INV_X1    g0311(.A(new_n492), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G97), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n318), .A2(new_n319), .A3(G244), .A4(new_n279), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n285), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n457), .A2(G257), .A3(new_n292), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n521), .A2(G190), .A3(new_n466), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n466), .A3(new_n522), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n511), .A2(new_n513), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n267), .A2(new_n500), .ZN(new_n527));
  AOI211_X1 g0327(.A(new_n508), .B(new_n505), .C1(new_n506), .C2(G107), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n513), .C1(new_n528), .C2(new_n383), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n521), .A2(new_n466), .A3(new_n522), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n438), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n303), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n490), .A2(new_n493), .A3(new_n497), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n460), .A2(new_n295), .A3(new_n466), .ZN(new_n536));
  INV_X1    g0336(.A(new_n466), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n459), .A2(KEYINPUT90), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n470), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(G200), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n498), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT83), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT19), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n546), .A3(new_n369), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n217), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n342), .A2(new_n500), .A3(new_n249), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n217), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n278), .A2(new_n217), .A3(G68), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(new_n546), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n396), .B2(new_n500), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n264), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n390), .A2(new_n418), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n318), .A2(new_n319), .A3(G238), .A4(new_n279), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n318), .A2(new_n319), .A3(G244), .A4(G1698), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n253), .C2(new_n207), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n285), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n292), .B(G250), .C1(G1), .C2(new_n455), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n456), .A2(G274), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n492), .A2(KEYINPUT85), .A3(new_n342), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT85), .B1(new_n492), .B2(new_n342), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n558), .A2(new_n559), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n566), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G190), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n557), .A2(new_n264), .B1(new_n390), .B2(new_n418), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n567), .A4(new_n570), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n318), .A2(new_n319), .A3(G257), .A4(new_n279), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n318), .A2(new_n319), .A3(G264), .A4(G1698), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n278), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n285), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n457), .A2(G270), .A3(new_n292), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n466), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n390), .A2(new_n207), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n207), .B1(new_n216), .B2(G33), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n383), .A2(new_n384), .A3(new_n386), .A4(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n263), .A2(new_n229), .B1(G20), .B2(new_n207), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n519), .B(new_n217), .C1(G33), .C2(new_n500), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(G169), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n593), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n585), .A2(KEYINPUT21), .A3(G169), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n583), .A2(G179), .A3(new_n466), .A4(new_n584), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n418), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n512), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n576), .A2(new_n605), .B1(new_n303), .B2(new_n566), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n574), .A2(new_n438), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n585), .A2(G200), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n609), .B(new_n598), .C1(new_n295), .C2(new_n585), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n578), .A2(new_n603), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n542), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n445), .A2(new_n612), .ZN(G372));
  NOR2_X1   g0413(.A1(new_n597), .A2(new_n602), .ZN(new_n614));
  INV_X1    g0414(.A(new_n601), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n467), .B1(new_n539), .B2(G179), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n535), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n571), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n606), .A2(new_n607), .B1(new_n618), .B2(new_n575), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n617), .A2(new_n541), .A3(new_n534), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n533), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n578), .A2(new_n621), .A3(new_n608), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n533), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT91), .A4(new_n532), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n619), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n620), .A2(new_n623), .A3(new_n608), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n445), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n414), .A2(new_n440), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n354), .A3(new_n401), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n340), .A2(new_n351), .ZN(new_n634));
  INV_X1    g0434(.A(new_n357), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT92), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT92), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n358), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(KEYINPUT18), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n358), .A2(new_n638), .ZN(new_n641));
  AOI211_X1 g0441(.A(KEYINPUT92), .B(new_n357), .C1(new_n340), .C2(new_n351), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n360), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n302), .B1(new_n633), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT93), .B1(new_n645), .B2(new_n306), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n645), .A2(KEYINPUT93), .A3(new_n306), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n631), .B1(new_n647), .B2(new_n648), .ZN(G369));
  AND2_X1   g0449(.A1(new_n498), .A2(new_n541), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT94), .B(KEYINPUT27), .Z(new_n651));
  NOR3_X1   g0451(.A1(new_n223), .A2(G1), .A3(G20), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n223), .A2(G20), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n216), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n650), .B1(new_n535), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n498), .B2(new_n659), .ZN(new_n661));
  INV_X1    g0461(.A(new_n603), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n598), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n603), .A2(new_n610), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n603), .A2(new_n658), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n650), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n498), .B2(new_n658), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  NOR2_X1   g0474(.A1(new_n224), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n551), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n228), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n617), .A2(new_n541), .A3(new_n619), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT97), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n526), .A2(new_n682), .A3(new_n533), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n526), .B2(new_n533), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI221_X1 g0485(.A(new_n608), .B1(KEYINPUT26), .B2(new_n622), .C1(new_n681), .C2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n628), .B1(new_n627), .B2(new_n619), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT29), .B(new_n659), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n630), .A2(new_n659), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n524), .A2(new_n566), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n538), .A2(new_n470), .ZN(new_n694));
  INV_X1    g0494(.A(new_n600), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT30), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n693), .A2(new_n694), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n530), .B1(new_n694), .B2(new_n466), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n566), .B(new_n585), .C1(new_n701), .C2(KEYINPUT95), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n473), .A2(KEYINPUT95), .A3(new_n524), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n438), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n612), .B2(new_n659), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT96), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n700), .B(new_n710), .C1(new_n702), .C2(new_n704), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n709), .A2(new_n658), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n692), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n680), .B1(new_n715), .B2(G1), .ZN(G364));
  XNOR2_X1  g0516(.A(new_n654), .B(KEYINPUT98), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n216), .B1(new_n717), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n675), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n668), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n666), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n229), .B1(G20), .B2(new_n303), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n217), .A2(new_n295), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n438), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n295), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n728), .A2(G58), .B1(G50), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n217), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n281), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT100), .Z(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G159), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT101), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT32), .ZN(new_n741));
  INV_X1    g0541(.A(new_n278), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n438), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n725), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n342), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n729), .A2(G190), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n742), .B(new_n745), .C1(G68), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n732), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n249), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n217), .B1(new_n736), .B2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(G97), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n735), .A2(new_n741), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G294), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n278), .B1(new_n730), .B2(G326), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n581), .B2(new_n744), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n756), .B(new_n758), .C1(new_n746), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  INV_X1    g0561(.A(G329), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n733), .A2(new_n761), .B1(new_n737), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n749), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(G283), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n760), .B(new_n765), .C1(new_n766), .C2(new_n727), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n724), .B1(new_n754), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n224), .A2(new_n278), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n228), .A2(G45), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n246), .C2(new_n455), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n225), .A2(G355), .A3(new_n278), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(G116), .C2(new_n225), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT99), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n723), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n768), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n720), .C1(new_n666), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n722), .A2(new_n781), .ZN(G396));
  NOR2_X1   g0582(.A1(new_n440), .A2(new_n658), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n426), .A2(new_n658), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n443), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n440), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n689), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n630), .A2(new_n659), .A3(new_n786), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n714), .B(new_n790), .Z(new_n791));
  INV_X1    g0591(.A(new_n720), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n749), .A2(new_n212), .ZN(new_n794));
  INV_X1    g0594(.A(G58), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n278), .B1(new_n751), .B2(new_n795), .C1(new_n744), .C2(new_n202), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n746), .A2(G150), .B1(new_n730), .B2(G137), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT103), .Z(new_n798));
  NAND2_X1  g0598(.A1(new_n728), .A2(G143), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n310), .C2(new_n733), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT104), .Z(new_n801));
  AOI211_X1 g0601(.A(new_n794), .B(new_n796), .C1(new_n801), .C2(KEYINPUT34), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(KEYINPUT34), .B2(new_n801), .C1(new_n803), .C2(new_n737), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n742), .B1(new_n751), .B2(new_n500), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  INV_X1    g0606(.A(new_n746), .ZN(new_n807));
  INV_X1    g0607(.A(new_n730), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n581), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n805), .B(new_n809), .C1(G311), .C2(new_n738), .ZN(new_n810));
  INV_X1    g0610(.A(new_n744), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G107), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n764), .A2(G87), .ZN(new_n813));
  INV_X1    g0613(.A(new_n733), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G294), .A2(new_n728), .B1(new_n814), .B2(G116), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n724), .B1(new_n804), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n723), .A2(new_n774), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n281), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n720), .C1(new_n776), .C2(new_n786), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n793), .A2(new_n820), .ZN(G384));
  INV_X1    g0621(.A(KEYINPUT40), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n330), .A2(new_n264), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n327), .A2(G68), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT79), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n327), .A2(KEYINPUT79), .A3(G68), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT16), .B1(new_n828), .B2(new_n312), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n351), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n656), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n362), .ZN(new_n834));
  INV_X1    g0634(.A(new_n363), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n636), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT17), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n353), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n833), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n311), .B1(new_n826), .B2(new_n827), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n383), .B1(new_n842), .B2(KEYINPUT16), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n312), .B1(new_n328), .B2(new_n329), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n331), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n350), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n353), .B1(new_n846), .B2(new_n656), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n357), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n634), .A2(new_n831), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n636), .A2(new_n850), .A3(new_n851), .A4(new_n353), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n841), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n854));
  INV_X1    g0654(.A(new_n850), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n640), .A2(new_n643), .A3(new_n354), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n637), .A2(new_n639), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(new_n353), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n855), .A2(new_n856), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n658), .A4(new_n711), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n708), .B2(new_n712), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n414), .A2(new_n401), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n412), .A2(new_n658), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n414), .A2(new_n401), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n863), .A2(new_n786), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n822), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n832), .B1(new_n365), .B2(new_n354), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n850), .A2(new_n851), .A3(new_n353), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n830), .A2(new_n635), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n832), .A2(new_n876), .A3(new_n353), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n636), .A2(new_n875), .B1(new_n877), .B2(KEYINPUT37), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n873), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT107), .A3(new_n854), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n841), .A2(new_n853), .A3(new_n881), .A4(KEYINPUT38), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n870), .A2(new_n880), .A3(new_n822), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n872), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n445), .A2(new_n863), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(G330), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n879), .A2(KEYINPUT107), .A3(new_n854), .ZN(new_n888));
  INV_X1    g0688(.A(new_n882), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n414), .A2(new_n658), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n861), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n783), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n789), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT106), .B1(new_n789), .B2(new_n895), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(new_n869), .A3(new_n880), .A4(new_n882), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n644), .A2(new_n831), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n887), .B(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n445), .A2(new_n691), .A3(new_n688), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n648), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n646), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n905), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n216), .B2(new_n717), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n503), .A2(new_n504), .ZN(new_n912));
  OAI211_X1 g0712(.A(G20), .B(new_n289), .C1(new_n912), .C2(KEYINPUT35), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n207), .B(new_n913), .C1(KEYINPUT35), .C2(new_n912), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT105), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI21_X1  g0716(.A(G77), .B1(new_n795), .B2(new_n212), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n917), .A2(new_n228), .B1(G50), .B2(new_n212), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n223), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n916), .A3(new_n919), .ZN(G367));
  INV_X1    g0720(.A(new_n769), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n778), .B1(new_n225), .B2(new_n418), .C1(new_n241), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n748), .ZN(new_n923));
  AOI22_X1  g0723(.A1(G97), .A2(new_n923), .B1(new_n814), .B2(G283), .ZN(new_n924));
  INV_X1    g0724(.A(G317), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n925), .B2(new_n737), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n730), .A2(G311), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n752), .A2(G107), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT46), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n744), .B2(new_n207), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n742), .B1(new_n807), .B2(new_n755), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n926), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n728), .A2(G303), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n738), .A2(G137), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n202), .B2(new_n733), .C1(new_n260), .C2(new_n727), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n278), .B1(new_n744), .B2(new_n795), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n746), .A2(G159), .B1(new_n730), .B2(G143), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n212), .B2(new_n751), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n923), .A2(G77), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n934), .A2(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT47), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n792), .B1(new_n944), .B2(new_n723), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n576), .A2(new_n570), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n658), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n619), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n608), .B2(new_n947), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n922), .B(new_n945), .C1(new_n949), .C2(new_n780), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT108), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n529), .A2(new_n658), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n683), .B2(new_n684), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n621), .A2(new_n658), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n673), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT44), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n673), .A2(new_n955), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n669), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n672), .B1(new_n661), .B2(new_n671), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n668), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n715), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n715), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n675), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n719), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n672), .A2(new_n953), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT42), .Z(new_n972));
  OR2_X1    g0772(.A1(new_n953), .A2(new_n498), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n658), .B1(new_n973), .B2(new_n533), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n970), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n955), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n670), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n951), .B1(new_n969), .B2(new_n980), .ZN(G387));
  NAND2_X1  g0781(.A1(new_n963), .A2(new_n719), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n738), .A2(G326), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n814), .A2(G303), .B1(G322), .B2(new_n730), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n761), .B2(new_n807), .C1(new_n925), .C2(new_n727), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT48), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n806), .B2(new_n751), .C1(new_n755), .C2(new_n744), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT49), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n278), .B(new_n983), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n988), .B2(new_n987), .C1(new_n207), .C2(new_n748), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n733), .A2(new_n212), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n752), .A2(new_n604), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n807), .B2(new_n255), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n742), .B(new_n993), .C1(G159), .C2(new_n730), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n811), .A2(G77), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n202), .B2(new_n727), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n764), .B2(G97), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(new_n260), .C2(new_n737), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n990), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n677), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n225), .A3(new_n278), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(G68), .B2(G77), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n256), .A2(new_n202), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n455), .C1(new_n1003), .C2(KEYINPUT50), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n769), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT109), .Z(new_n1007));
  NOR2_X1   g0807(.A1(new_n238), .A2(new_n455), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1001), .B1(G107), .B2(new_n225), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n999), .A2(new_n723), .B1(new_n778), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n720), .C1(new_n661), .C2(new_n780), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n675), .B1(new_n963), .B2(new_n715), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n982), .B(new_n1011), .C1(new_n965), .C2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT110), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(G393));
  INV_X1    g0815(.A(new_n961), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n964), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n966), .A2(new_n1017), .A3(new_n675), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n961), .A2(new_n719), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n778), .B1(new_n500), .B2(new_n225), .C1(new_n251), .C2(new_n921), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n751), .A2(new_n281), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n278), .B1(new_n733), .B2(new_n255), .C1(new_n212), .C2(new_n744), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G50), .C2(new_n746), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n808), .A2(new_n260), .B1(new_n727), .B2(new_n310), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n738), .A2(G143), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n813), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n742), .B1(new_n737), .B2(new_n766), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n807), .A2(new_n581), .B1(new_n751), .B2(new_n207), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G294), .C2(new_n814), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n808), .A2(new_n925), .B1(new_n727), .B2(new_n761), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(new_n249), .C2(new_n749), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n744), .A2(new_n806), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n792), .B1(new_n1036), .B2(new_n723), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1020), .B(new_n1037), .C1(new_n976), .C2(new_n780), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1018), .A2(new_n1019), .A3(new_n1038), .ZN(G390));
  NAND3_X1  g0839(.A1(new_n445), .A2(G330), .A3(new_n863), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n870), .A2(G330), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n869), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n714), .B2(new_n787), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1041), .A2(new_n1043), .B1(new_n899), .B2(new_n897), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n863), .A2(G330), .A3(new_n786), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n785), .A2(new_n440), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n659), .B(new_n1047), .C1(new_n686), .C2(new_n687), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1048), .A2(new_n895), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n713), .A2(new_n869), .A3(G330), .A4(new_n786), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n909), .B(new_n1040), .C1(new_n1044), .C2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n869), .B1(new_n896), .B2(new_n898), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n891), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n892), .B1(new_n880), .B2(new_n882), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n856), .A2(new_n855), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n859), .A2(new_n852), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n873), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT39), .B1(new_n1061), .B2(new_n854), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1056), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n861), .B(new_n1055), .C1(new_n1049), .C2(new_n1042), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1050), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1041), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1053), .B(new_n1066), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n906), .B(new_n1040), .C1(new_n647), .C2(new_n648), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n900), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1070), .B1(new_n1072), .B2(new_n1051), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1068), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1069), .A2(new_n1076), .A3(new_n675), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n775), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n738), .A2(G125), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1079), .B1(new_n803), .B2(new_n727), .C1(new_n733), .C2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n742), .B(new_n1082), .C1(G137), .C2(new_n746), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n730), .A2(G128), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n811), .A2(G150), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1084), .B1(new_n310), .B2(new_n751), .C1(new_n1085), .C2(KEYINPUT53), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(KEYINPUT53), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1087), .C1(new_n202), .C2(new_n748), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n727), .A2(new_n207), .B1(new_n733), .B2(new_n500), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n794), .A2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n807), .A2(new_n249), .B1(new_n808), .B2(new_n806), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1091), .A2(new_n745), .A3(new_n278), .A4(new_n1021), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n755), .C2(new_n737), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n724), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n255), .B2(new_n818), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1078), .A2(new_n720), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n719), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1077), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT112), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT112), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1077), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(G378));
  NOR2_X1   g0903(.A1(new_n273), .A2(new_n656), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n307), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1105), .B(new_n1106), .Z(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G330), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n872), .B2(new_n883), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n904), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n883), .ZN(new_n1114));
  OAI21_X1  g0914(.A(G330), .B1(new_n1114), .B2(new_n871), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n902), .B1(new_n1116), .B2(new_n891), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n901), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1070), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1076), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n904), .A2(new_n1112), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n901), .A3(new_n1115), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1119), .A2(new_n1121), .A3(KEYINPUT57), .A4(new_n1124), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n675), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1081), .A2(new_n744), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(KEYINPUT114), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G150), .B2(new_n752), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1130), .A2(KEYINPUT114), .B1(G137), .B2(new_n814), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n728), .A2(G128), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n746), .A2(G132), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G125), .B2(new_n730), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT59), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n923), .A2(G159), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G33), .B1(new_n738), .B2(G124), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n733), .A2(new_n418), .B1(new_n737), .B2(new_n806), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n728), .A2(KEYINPUT113), .A3(G107), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT113), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n727), .B2(new_n249), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n746), .A2(G97), .B1(new_n730), .B2(G116), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n278), .B1(new_n752), .B2(G68), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n995), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n748), .A2(new_n795), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT58), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n1143), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT58), .B1(new_n1153), .B2(new_n287), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1157));
  AOI21_X1  g0957(.A(G50), .B1(new_n1157), .B2(new_n287), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(new_n723), .B1(new_n202), .B2(new_n818), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1109), .B2(new_n776), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(new_n792), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1122), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1109), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1162), .B1(new_n1165), .B2(new_n719), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1129), .A2(new_n1166), .ZN(G375));
  NOR2_X1   g0967(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1168), .A2(KEYINPUT117), .A3(new_n1070), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT117), .B1(new_n1168), .B2(new_n1070), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n968), .B(new_n1053), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1168), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n818), .A2(new_n212), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n869), .A2(G13), .A3(G33), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n742), .B1(new_n749), .B2(new_n281), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT119), .Z(new_n1176));
  OAI22_X1  g0976(.A1(new_n744), .A2(new_n500), .B1(new_n737), .B2(new_n581), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT120), .Z(new_n1178));
  AND3_X1   g0978(.A1(new_n1176), .A2(new_n992), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n746), .A2(G116), .B1(new_n730), .B2(G294), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n249), .B2(new_n733), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n806), .C2(new_n727), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT121), .Z(new_n1184));
  OAI22_X1  g0984(.A1(new_n744), .A2(new_n310), .B1(new_n733), .B2(new_n260), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G137), .B2(new_n728), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n738), .A2(G128), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n742), .B1(new_n746), .B2(new_n1080), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n808), .A2(new_n803), .B1(new_n751), .B2(new_n202), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(new_n1152), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n724), .B1(new_n1184), .B2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1174), .A2(new_n792), .A3(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1172), .A2(new_n719), .B1(new_n1173), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1171), .A2(new_n1194), .ZN(G381));
  XNOR2_X1  g0995(.A(G375), .B(KEYINPUT123), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1099), .ZN(new_n1197));
  INV_X1    g0997(.A(G381), .ZN(new_n1198));
  INV_X1    g0998(.A(G396), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1014), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT122), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1202), .A2(G387), .A3(G390), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1203), .ZN(G407));
  NAND3_X1  g1004(.A1(new_n1196), .A2(new_n657), .A3(new_n1197), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(G407), .A2(G213), .A3(new_n1205), .ZN(G409));
  AND2_X1   g1006(.A1(new_n657), .A2(G213), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT124), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1119), .A2(new_n1209), .A3(new_n1124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1210), .A3(new_n719), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1162), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1165), .A2(new_n968), .A3(new_n1121), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1197), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1129), .A2(G378), .A3(new_n1166), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1207), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1053), .A2(KEYINPUT60), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1070), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n675), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(G384), .A3(new_n1194), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G384), .B1(new_n1221), .B2(new_n1194), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G2897), .B(new_n1207), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1224), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1207), .A2(G2897), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1222), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT63), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1222), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1217), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G387), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G390), .B(new_n951), .C1(new_n969), .C2(new_n980), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1014), .B(G396), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1235), .A2(G387), .A3(KEYINPUT126), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1235), .A2(G387), .A3(KEYINPUT125), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n1240), .A3(new_n1237), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1207), .B(new_n1231), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(KEYINPUT63), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1234), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1217), .A2(new_n1253), .A3(new_n1232), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1217), .B2(new_n1232), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1248), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1252), .B1(new_n1257), .B2(new_n1258), .ZN(G405));
  AOI21_X1  g1059(.A(new_n1099), .B1(new_n1129), .B2(new_n1166), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT127), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1231), .B1(new_n1261), .B2(new_n1216), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1197), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT127), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1266));
  AND4_X1   g1066(.A1(new_n1216), .A2(new_n1264), .A3(new_n1231), .A4(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1248), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1216), .A3(new_n1231), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1216), .A3(new_n1266), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1232), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1271), .A3(new_n1258), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(G402));
endmodule


