//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n190), .B(KEYINPUT1), .C1(new_n187), .C2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G128), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n187), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n194), .A3(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT65), .A3(new_n198), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n192), .A2(new_n196), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n196), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT80), .B1(new_n211), .B2(new_n205), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G125), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n216), .A2(G224), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n206), .A2(new_n212), .A3(new_n215), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n201), .A2(new_n203), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n191), .A2(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n190), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n196), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  MUX2_X1   g039(.A(new_n211), .B(new_n225), .S(new_n205), .Z(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n226), .B2(new_n219), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n228), .B(KEYINPUT8), .Z(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G116), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(G113), .B(new_n232), .C1(new_n234), .C2(new_n230), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n239), .B2(G107), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  INV_X1    g055(.A(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G104), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(G107), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n239), .A2(G107), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(G104), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n235), .A2(new_n238), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n246), .A2(new_n249), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n235), .A3(new_n238), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(KEYINPUT81), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n252), .A2(KEYINPUT81), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n229), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n227), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n243), .A3(new_n245), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n234), .A2(new_n236), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n238), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n262), .A3(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT79), .A4(new_n263), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n228), .A3(new_n252), .A4(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n256), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n252), .A3(new_n267), .ZN(new_n270));
  INV_X1    g084(.A(new_n228), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT6), .A3(new_n268), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n206), .A2(new_n212), .A3(new_n215), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(new_n217), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n269), .A2(new_n280), .A3(new_n278), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G214), .B1(G237), .B2(G902), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT78), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT9), .B(G234), .ZN(new_n288));
  OAI21_X1  g102(.A(G221), .B1(new_n288), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G110), .B(G140), .ZN(new_n294));
  INV_X1    g108(.A(G227), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n259), .A2(new_n263), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n211), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n246), .A2(new_n249), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n225), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n188), .A2(G128), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n196), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT65), .B1(new_n202), .B2(new_n198), .ZN(new_n308));
  AND4_X1   g122(.A1(KEYINPUT65), .A2(new_n198), .A3(new_n194), .A4(new_n195), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n310), .B2(new_n251), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n188), .A2(G128), .B1(new_n194), .B2(new_n195), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n201), .B2(new_n203), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(KEYINPUT76), .A3(new_n300), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n301), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n313), .B2(new_n300), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n305), .A3(new_n251), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT77), .A3(new_n301), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n304), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT64), .B1(new_n323), .B2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT64), .B(new_n326), .C1(new_n323), .C2(G137), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n331), .A3(new_n327), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n297), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n299), .A2(new_n303), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n320), .B2(new_n301), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n316), .B(KEYINPUT10), .C1(new_n318), .C2(new_n319), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n333), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n334), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n311), .A2(new_n314), .B1(new_n225), .B2(new_n251), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT12), .A3(new_n333), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n318), .A2(new_n319), .B1(new_n204), .B2(new_n300), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n335), .A2(new_n340), .B1(new_n348), .B2(new_n297), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n293), .B1(new_n349), .B2(G469), .ZN(new_n350));
  INV_X1    g164(.A(new_n297), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n340), .B2(new_n341), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n341), .A2(new_n347), .A3(new_n351), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n291), .B(new_n292), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n290), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n287), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G125), .B(G140), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n358));
  OR3_X1    g172(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(G146), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n216), .A3(G214), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n187), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(G214), .C1(KEYINPUT83), .C2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G131), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n331), .A3(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n331), .B1(new_n366), .B2(new_n368), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n374), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT86), .B1(new_n374), .B2(KEYINPUT17), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n362), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n357), .B(new_n193), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n369), .A2(KEYINPUT84), .A3(new_n378), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT84), .B1(new_n369), .B2(new_n378), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n379), .B(new_n380), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G113), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n239), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n377), .A2(new_n384), .ZN(new_n389));
  INV_X1    g203(.A(new_n386), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT87), .B(new_n386), .C1(new_n377), .C2(new_n384), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n292), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n370), .A2(new_n372), .ZN(new_n395));
  INV_X1    g209(.A(new_n360), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n357), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n193), .C1(new_n357), .C2(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n384), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n390), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n387), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n411), .A3(new_n406), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n394), .A2(G475), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT15), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G478), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n187), .A2(G128), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n197), .A2(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n323), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n418), .A3(G134), .ZN(new_n421));
  OR2_X1    g235(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n418), .A3(G134), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n422), .A2(new_n423), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(G134), .A3(new_n417), .A4(new_n418), .ZN(new_n427));
  INV_X1    g241(.A(G122), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT88), .B1(new_n428), .B2(G116), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  INV_X1    g244(.A(G116), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(G116), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n433), .A2(new_n242), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n242), .B1(new_n433), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n425), .B(new_n427), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n420), .A2(new_n421), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n433), .A2(KEYINPUT14), .B1(G116), .B2(new_n428), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n242), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n437), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G217), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n288), .A2(new_n445), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n441), .A2(new_n442), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n439), .B1(new_n449), .B2(new_n242), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n437), .A3(new_n446), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n416), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n416), .B1(new_n452), .B2(new_n453), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(G234), .A2(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(G952), .A3(new_n216), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT91), .Z(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(G898), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT92), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n461), .A2(G902), .A3(G953), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n414), .A2(new_n460), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n356), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n323), .A2(G137), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n323), .A2(G137), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n332), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n225), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(KEYINPUT11), .B2(new_n324), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n331), .B1(new_n477), .B2(new_n327), .ZN(new_n478));
  INV_X1    g292(.A(new_n332), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n211), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n261), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n476), .B2(new_n480), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT28), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n367), .A2(G210), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT26), .B(G101), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n476), .A2(new_n480), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n481), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n333), .A2(new_n211), .B1(new_n475), .B2(new_n225), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(KEYINPUT30), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n476), .A2(new_n480), .A3(new_n498), .A4(KEYINPUT30), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n491), .B1(new_n503), .B2(new_n482), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n292), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n485), .A2(KEYINPUT29), .A3(new_n487), .A4(new_n491), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT28), .B1(new_n499), .B2(new_n481), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n332), .A2(new_n474), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n204), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n213), .B1(new_n330), .B2(new_n332), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n261), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n482), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n513), .B2(KEYINPUT28), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT29), .A4(new_n491), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G472), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n491), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n503), .A2(new_n520), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n521), .A2(KEYINPUT31), .B1(new_n514), .B2(new_n491), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n476), .A2(new_n480), .A3(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT67), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n501), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n519), .B1(new_n526), .B2(new_n497), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT31), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n522), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n518), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n485), .A2(new_n487), .ZN(new_n538));
  INV_X1    g352(.A(new_n491), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n527), .A2(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT68), .B1(new_n521), .B2(KEYINPUT31), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n527), .A2(new_n523), .A3(new_n528), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT32), .B1(new_n543), .B2(new_n532), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT70), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n445), .B1(G234), .B2(new_n292), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n357), .A2(new_n193), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n231), .A2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n197), .A2(G119), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT71), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  INV_X1    g368(.A(new_n549), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n548), .B(new_n554), .C1(new_n555), .C2(KEYINPUT23), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n396), .B(new_n547), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(G110), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n560), .C1(new_n360), .C2(new_n361), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT22), .B(G137), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n558), .A2(new_n561), .A3(new_n565), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n567), .A2(new_n292), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT72), .B1(KEYINPUT73), .B2(KEYINPUT25), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n546), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n567), .A2(new_n572), .A3(new_n292), .A4(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT25), .B1(new_n573), .B2(KEYINPUT73), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n546), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n292), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n567), .A2(new_n568), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n483), .B1(new_n526), .B2(new_n497), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n493), .B(new_n492), .C1(new_n582), .C2(new_n491), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(new_n292), .A3(new_n507), .A4(new_n516), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n543), .A2(new_n535), .B1(new_n584), .B2(G472), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n534), .B1(new_n531), .B2(new_n533), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n545), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT75), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n545), .A2(new_n588), .A3(new_n591), .A4(new_n581), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n471), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n244), .ZN(G3));
  NOR2_X1   g408(.A1(new_n531), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n531), .A2(new_n533), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n581), .A3(new_n355), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n448), .A2(new_n451), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n448), .A2(KEYINPUT33), .A3(new_n451), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n607));
  OAI21_X1  g421(.A(G478), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n292), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n452), .B2(new_n609), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n413), .ZN(new_n613));
  INV_X1    g427(.A(new_n285), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n282), .B2(new_n283), .ZN(new_n615));
  INV_X1    g429(.A(new_n469), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n600), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  XNOR2_X1  g434(.A(new_n407), .B(new_n409), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n394), .A2(G475), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n615), .A2(new_n624), .A3(new_n616), .A4(new_n460), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n600), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  INV_X1    g443(.A(new_n456), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n454), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n458), .B1(new_n631), .B2(new_n416), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n562), .A2(KEYINPUT96), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n558), .A2(new_n635), .A3(new_n561), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n634), .B1(new_n633), .B2(new_n636), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n578), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n571), .B2(new_n574), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n632), .A2(new_n413), .A3(new_n640), .A4(new_n616), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n597), .A2(new_n598), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n356), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(new_n293), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n335), .A2(new_n340), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n348), .A2(new_n297), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(G469), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n354), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n289), .A2(new_n650), .A3(new_n615), .A4(new_n640), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n216), .A2(G900), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(G902), .A3(new_n461), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT97), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n463), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n623), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n460), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n651), .A2(new_n545), .A3(new_n588), .A4(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NAND2_X1  g478(.A1(new_n282), .A2(new_n283), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n460), .A2(new_n285), .ZN(new_n668));
  OR4_X1    g482(.A1(new_n413), .A2(new_n667), .A3(new_n640), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n655), .B(KEYINPUT39), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n355), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT40), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n543), .A2(new_n535), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n582), .A2(new_n539), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n292), .B1(new_n513), .B2(new_n491), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n586), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT99), .ZN(new_n680));
  OR3_X1    g494(.A1(new_n669), .A2(new_n672), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  INV_X1    g496(.A(new_n612), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n414), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n656), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n651), .A2(new_n545), .A3(new_n588), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NOR3_X1   g501(.A1(new_n537), .A2(new_n544), .A3(KEYINPUT70), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n587), .B1(new_n585), .B2(new_n586), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n292), .B1(new_n352), .B2(new_n353), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n289), .A3(new_n354), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n617), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n690), .A2(KEYINPUT100), .A3(new_n581), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n617), .A2(new_n693), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n589), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NOR2_X1   g515(.A1(new_n625), .A2(new_n693), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n545), .A3(new_n581), .A4(new_n588), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  INV_X1    g518(.A(new_n615), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n693), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n641), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n545), .A2(new_n706), .A3(new_n588), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  XOR2_X1   g523(.A(new_n532), .B(KEYINPUT101), .Z(new_n710));
  NOR2_X1   g524(.A1(new_n527), .A2(new_n528), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n522), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n581), .B(new_n712), .C1(new_n595), .C2(new_n596), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n284), .A2(new_n668), .A3(new_n413), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n693), .A2(new_n469), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  OAI211_X1 g532(.A(new_n640), .B(new_n712), .C1(new_n595), .C2(new_n596), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n685), .A3(new_n706), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n650), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n665), .A2(new_n290), .A3(new_n614), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n350), .A2(KEYINPUT102), .A3(new_n354), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n589), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n685), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n685), .A2(new_n724), .A3(new_n725), .A4(new_n726), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n585), .A2(new_n586), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n581), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT42), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n685), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n589), .A2(new_n737), .A3(KEYINPUT42), .A4(new_n727), .ZN(new_n738));
  INV_X1    g552(.A(new_n735), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT103), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n331), .ZN(G33));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n728), .B2(new_n659), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n589), .A2(new_n658), .A3(new_n727), .A4(KEYINPUT104), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  OR2_X1    g561(.A1(new_n349), .A2(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n349), .A2(KEYINPUT45), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(G469), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n646), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n646), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n354), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(new_n289), .A3(new_n670), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n683), .A2(new_n413), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n414), .A2(KEYINPUT43), .A3(new_n612), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n640), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n599), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n665), .A2(new_n614), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n761), .B2(KEYINPUT44), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n756), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(G137), .Z(G39));
  NOR4_X1   g581(.A1(new_n690), .A2(new_n581), .A3(new_n737), .A4(new_n764), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT105), .Z(new_n769));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n289), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT106), .B(G140), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G42));
  NAND2_X1  g589(.A1(new_n759), .A2(new_n758), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n713), .A3(new_n463), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n706), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT115), .Z(new_n779));
  NAND2_X1  g593(.A1(new_n692), .A2(new_n354), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n464), .A3(new_n725), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n680), .A2(new_n581), .A3(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(G952), .B(new_n216), .C1(new_n784), .C2(new_n684), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n782), .A2(new_n734), .A3(new_n776), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT48), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n779), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n666), .A2(new_n285), .A3(new_n693), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT50), .Z(new_n791));
  NAND4_X1  g605(.A1(new_n783), .A2(new_n720), .A3(new_n758), .A4(new_n759), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n612), .A2(new_n413), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n791), .B(new_n792), .C1(new_n784), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n772), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n289), .B2(new_n780), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n777), .A2(new_n763), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n788), .B1(new_n798), .B2(KEYINPUT51), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT114), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT114), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n732), .A2(new_n719), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n632), .A2(new_n640), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n355), .A2(new_n657), .A3(new_n763), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n804), .B1(new_n690), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n744), .B2(new_n745), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT109), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n810), .B(new_n807), .C1(new_n744), .C2(new_n745), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n741), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n684), .B1(new_n414), .B2(new_n632), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n287), .A3(new_n616), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n643), .B1(new_n600), .B2(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n593), .A2(KEYINPUT108), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT108), .B1(new_n593), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n703), .A2(new_n717), .A3(new_n708), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n699), .A2(new_n819), .A3(KEYINPUT107), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT107), .B1(new_n699), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n655), .A2(new_n289), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n640), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n724), .A2(new_n726), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n724), .A2(new_n826), .A3(KEYINPUT110), .A4(new_n726), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n715), .B1(new_n544), .B2(new_n677), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT111), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n835), .B(new_n832), .C1(new_n829), .C2(new_n830), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n721), .A2(new_n686), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n823), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(KEYINPUT102), .A2(new_n354), .A3(new_n646), .A4(new_n649), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT102), .B1(new_n350), .B2(new_n354), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT110), .B1(new_n845), .B2(new_n826), .ZN(new_n846));
  INV_X1    g660(.A(new_n830), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n833), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n835), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n831), .A2(KEYINPUT111), .A3(new_n833), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n721), .A2(new_n686), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n661), .B2(new_n662), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n812), .A2(new_n818), .A3(new_n822), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n837), .A2(new_n841), .A3(new_n823), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n851), .B2(new_n853), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n818), .B(new_n822), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n809), .A2(new_n811), .ZN(new_n862));
  INV_X1    g676(.A(new_n741), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n857), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(KEYINPUT112), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n867), .A3(new_n857), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n699), .A2(new_n819), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n871), .A2(new_n857), .A3(new_n739), .A4(new_n738), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n862), .A2(new_n818), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n855), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n857), .C1(new_n861), .C2(new_n864), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n856), .B2(new_n857), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n870), .B(new_n876), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n803), .A2(new_n869), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n885));
  INV_X1    g699(.A(new_n286), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n581), .A2(new_n289), .A3(new_n886), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n884), .A2(new_n885), .A3(new_n757), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n680), .A2(new_n888), .A3(new_n667), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n875), .B1(new_n891), .B2(new_n878), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n292), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n273), .A2(new_n275), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n277), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  NOR2_X1   g711(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n216), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  XNOR2_X1  g716(.A(new_n293), .B(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n891), .B2(new_n878), .ZN(new_n905));
  OAI22_X1  g719(.A1(KEYINPUT117), .A2(new_n905), .B1(new_n892), .B2(new_n870), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(KEYINPUT117), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n352), .A2(new_n353), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n750), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT118), .B1(new_n893), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n913));
  AND4_X1   g727(.A1(KEYINPUT118), .A2(new_n913), .A3(G902), .A4(new_n911), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n901), .B1(new_n910), .B2(new_n915), .ZN(G54));
  INV_X1    g730(.A(new_n901), .ZN(new_n917));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(G902), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n405), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT120), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n913), .A2(G902), .A3(new_n405), .A4(new_n918), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT119), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(G60));
  XNOR2_X1  g740(.A(new_n610), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n869), .B2(new_n881), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n606), .A2(new_n607), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT121), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n917), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n906), .A2(new_n907), .ZN(new_n932));
  INV_X1    g746(.A(new_n927), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n892), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n637), .B2(new_n638), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n579), .B1(new_n892), .B2(new_n937), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n917), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n917), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n216), .B1(new_n466), .B2(G224), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n818), .A2(new_n822), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n216), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n895), .B1(G898), .B2(new_n216), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(G69));
  OAI21_X1  g764(.A(new_n526), .B1(KEYINPUT30), .B2(new_n499), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT122), .Z(new_n952));
  OAI21_X1  g766(.A(new_n400), .B1(new_n357), .B2(new_n399), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(new_n954));
  AOI21_X1  g768(.A(new_n766), .B1(new_n769), .B2(new_n772), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n863), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n756), .A2(new_n581), .A3(new_n733), .A4(new_n715), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n746), .A2(new_n853), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n216), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n652), .B(KEYINPUT124), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n954), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n681), .A2(new_n853), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT123), .Z(new_n965));
  OR2_X1    g779(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n590), .A2(new_n592), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n813), .A2(new_n763), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n355), .A3(new_n670), .A4(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n966), .A3(new_n969), .A4(new_n955), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n216), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n962), .B1(new_n971), .B2(new_n954), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n216), .B1(G227), .B2(G900), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(G72));
  NAND2_X1  g788(.A1(new_n582), .A2(new_n539), .ZN(new_n975));
  XOR2_X1   g789(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n976));
  NOR2_X1   g790(.A1(new_n596), .A2(new_n292), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n674), .A2(new_n978), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n868), .A2(new_n866), .A3(new_n975), .A4(new_n979), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n978), .B(KEYINPUT126), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n970), .B2(new_n947), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n674), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n956), .A2(new_n818), .A3(new_n822), .A4(new_n958), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n975), .B1(new_n985), .B2(new_n981), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(new_n901), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n986), .A2(new_n984), .A3(new_n901), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n980), .B(new_n983), .C1(new_n987), .C2(new_n988), .ZN(G57));
endmodule


