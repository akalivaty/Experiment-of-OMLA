//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT90), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT90), .A2(G952), .ZN(new_n189));
  AOI21_X1  g003(.A(G953), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G234), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT21), .B(G898), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(KEYINPUT91), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G902), .ZN(new_n198));
  INV_X1    g012(.A(G953), .ZN(new_n199));
  AOI211_X1 g013(.A(new_n198), .B(new_n199), .C1(G234), .C2(G237), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n194), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G210), .B1(G237), .B2(G902), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT76), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT76), .A4(G104), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n213), .B(KEYINPUT3), .C1(new_n204), .C2(G107), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(KEYINPUT3), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n214), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(new_n209), .A3(G104), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n210), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n222), .A2(new_n226), .A3(new_n227), .A4(new_n205), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n219), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(G116), .B(G119), .Z(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(G101), .C1(new_n212), .C2(new_n218), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G110), .B(G122), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT80), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n205), .A2(new_n216), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(G113), .C1(KEYINPUT5), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n235), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n241), .B(KEYINPUT8), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n244), .A2(new_n249), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n228), .A2(new_n243), .B1(new_n248), .B2(new_n235), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G128), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n262), .B(G146), .C1(new_n259), .C2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n256), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n256), .A2(new_n267), .ZN(new_n270));
  OAI21_X1  g084(.A(G125), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n199), .A2(G224), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n266), .A2(new_n271), .A3(new_n273), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OR3_X1    g092(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n274), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n251), .A2(new_n255), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n198), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n239), .A2(new_n250), .ZN(new_n284));
  INV_X1    g098(.A(new_n241), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n251), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n239), .A2(new_n241), .A3(new_n250), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n241), .B1(new_n239), .B2(new_n250), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n284), .A2(new_n290), .A3(new_n285), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n287), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n275), .A2(new_n276), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n283), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n281), .B1(new_n280), .B2(new_n198), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n203), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n286), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT81), .B1(new_n289), .B2(new_n290), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n304), .B2(new_n287), .ZN(new_n305));
  INV_X1    g119(.A(new_n203), .ZN(new_n306));
  NOR4_X1   g120(.A1(new_n305), .A2(new_n306), .A3(new_n299), .A4(new_n283), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n187), .B(new_n202), .C1(new_n301), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G478), .ZN(new_n312));
  INV_X1    g126(.A(G122), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n313), .B2(G116), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT14), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G122), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(G116), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n314), .A2(new_n317), .A3(KEYINPUT86), .A4(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n314), .A2(new_n318), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(G107), .C1(new_n320), .C2(KEYINPUT86), .ZN(new_n321));
  XNOR2_X1  g135(.A(G128), .B(G143), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(G122), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n325), .A3(new_n209), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n262), .A2(G128), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(G134), .C1(KEYINPUT13), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(new_n323), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT68), .B(G217), .Z(new_n337));
  XOR2_X1   g151(.A(KEYINPUT9), .B(G234), .Z(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n199), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n339), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n335), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT87), .A3(new_n342), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n336), .A2(KEYINPUT87), .A3(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n198), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n312), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n348), .A2(new_n312), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G475), .ZN(new_n352));
  NOR2_X1   g166(.A1(G237), .A2(G953), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(G143), .A3(G214), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G143), .B1(new_n353), .B2(G214), .ZN(new_n356));
  OAI21_X1  g170(.A(G131), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n354), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT17), .B(G131), .C1(new_n355), .C2(new_n356), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G125), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n265), .A2(G140), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n366), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n260), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n362), .A2(new_n363), .A3(new_n372), .A4(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT84), .B(G104), .Z(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n368), .B2(new_n369), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n260), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n373), .A2(G146), .ZN(new_n385));
  AND2_X1   g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n358), .A2(new_n354), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n386), .B1(new_n358), .B2(new_n354), .ZN(new_n388));
  OAI22_X1  g202(.A1(new_n384), .A2(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n376), .A2(new_n379), .A3(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n357), .A2(new_n360), .B1(new_n371), .B2(G146), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n373), .A2(KEYINPUT83), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT19), .B1(new_n392), .B2(new_n382), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n260), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n379), .B1(new_n396), .B2(new_n389), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n352), .B(new_n198), .C1(new_n390), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT20), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n376), .A2(new_n389), .A3(new_n379), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n384), .A2(new_n385), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n387), .A2(new_n388), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n401), .A2(new_n402), .B1(new_n391), .B2(new_n395), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n400), .B1(new_n403), .B2(new_n379), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n352), .A4(new_n198), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n400), .A2(KEYINPUT85), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n379), .B1(new_n376), .B2(new_n389), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n198), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(KEYINPUT85), .B(new_n379), .C1(new_n376), .C2(new_n389), .ZN(new_n411));
  OAI21_X1  g225(.A(G475), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n351), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n308), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G221), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n338), .B2(new_n198), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n228), .A2(KEYINPUT10), .A3(new_n264), .A4(new_n243), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n423), .A2(KEYINPUT11), .B1(new_n323), .B2(G137), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT11), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT64), .A4(G134), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n423), .A2(KEYINPUT11), .B1(new_n323), .B2(G137), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n428), .A2(new_n359), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n359), .B1(new_n428), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n422), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND4_X1   g246(.A1(KEYINPUT64), .A2(new_n425), .A3(new_n426), .A4(G134), .ZN(new_n433));
  AOI22_X1  g247(.A1(KEYINPUT64), .A2(new_n425), .B1(new_n426), .B2(G134), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G131), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n428), .A2(new_n359), .A3(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT65), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n228), .A2(new_n264), .A3(new_n243), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n269), .A2(new_n270), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n229), .A2(new_n444), .A3(new_n238), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n421), .A2(new_n439), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n440), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n264), .B1(new_n228), .B2(new_n243), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n431), .B2(new_n430), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n438), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n264), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n244), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n440), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n449), .A2(KEYINPUT12), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G140), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n199), .A2(G227), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n460), .B(new_n461), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n439), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n445), .A2(new_n442), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n419), .B(KEYINPUT77), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(new_n446), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n430), .A2(new_n431), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n454), .B2(new_n440), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n447), .A2(new_n448), .ZN(new_n472));
  OAI22_X1  g286(.A1(new_n471), .A2(new_n450), .B1(new_n472), .B2(new_n451), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n465), .A2(new_n466), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n439), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n463), .B1(new_n475), .B2(new_n458), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n476), .A3(new_n198), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT78), .A3(G469), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n467), .A2(new_n446), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n463), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n446), .A2(new_n456), .A3(new_n462), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n481), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G469), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n198), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT78), .B1(new_n477), .B2(G469), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n418), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n432), .A2(new_n438), .A3(new_n444), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n426), .A2(G134), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n323), .A2(G137), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n264), .A2(new_n437), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(KEYINPUT30), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n443), .B1(new_n436), .B2(new_n437), .ZN(new_n499));
  INV_X1    g313(.A(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(new_n236), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n236), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n353), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G101), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n236), .B1(new_n499), .B2(new_n500), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT28), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n492), .A2(new_n496), .ZN(new_n522));
  INV_X1    g336(.A(new_n504), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n517), .B1(new_n524), .B2(new_n505), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT29), .A3(new_n511), .A4(new_n518), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n527), .A3(new_n198), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G472), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n502), .A2(new_n505), .A3(new_n511), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT31), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n502), .A2(new_n532), .A3(new_n505), .A4(new_n511), .ZN(new_n533));
  INV_X1    g347(.A(new_n518), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n517), .B1(new_n505), .B2(new_n514), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n512), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(KEYINPUT32), .A3(new_n538), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n529), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n337), .B1(new_n191), .B2(G902), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT69), .Z(new_n545));
  NAND3_X1  g359(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT72), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT22), .B(G137), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n372), .A2(new_n375), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT71), .B1(new_n246), .B2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n259), .A2(G119), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT71), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n552), .B(new_n555), .C1(G119), .C2(new_n259), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT70), .B1(new_n246), .B2(G128), .ZN(new_n558));
  MUX2_X1   g372(.A(KEYINPUT70), .B(new_n558), .S(new_n553), .Z(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n550), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n559), .A2(new_n560), .B1(new_n556), .B2(G110), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n385), .B1(new_n371), .B2(G146), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n549), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n565), .A3(new_n549), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT25), .B1(new_n569), .B2(new_n198), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n562), .A2(new_n565), .A3(new_n549), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT25), .B(new_n198), .C1(new_n571), .C2(new_n566), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n545), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n544), .A2(new_n198), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n543), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n416), .A2(new_n491), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT92), .B(G101), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G3));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n343), .A2(new_n344), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n342), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n327), .A2(new_n335), .A3(KEYINPUT93), .A4(new_n341), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n340), .A3(KEYINPUT33), .A4(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(G478), .A3(new_n198), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT94), .B(G478), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n345), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n407), .A2(new_n412), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n308), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n488), .A2(new_n490), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n578), .A2(new_n418), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n537), .A2(new_n198), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n539), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  OAI21_X1  g418(.A(new_n414), .B1(new_n349), .B2(new_n350), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n308), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n606), .A2(new_n596), .A3(new_n597), .A4(new_n601), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(new_n209), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n607), .B(new_n609), .ZN(G9));
  INV_X1    g424(.A(new_n545), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT25), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n571), .A2(new_n566), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(G902), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(new_n572), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n562), .A2(new_n565), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n576), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT96), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n574), .A2(new_n622), .A3(new_n619), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n416), .A2(new_n491), .A3(new_n601), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G110), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  INV_X1    g443(.A(new_n418), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n478), .A2(new_n487), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n543), .B(new_n630), .C1(new_n631), .C2(new_n489), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n200), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n634), .A2(new_n193), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n605), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n625), .B(new_n187), .C1(new_n301), .C2(new_n307), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n259), .ZN(G30));
  XOR2_X1   g454(.A(new_n635), .B(KEYINPUT39), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n491), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT40), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n301), .A2(new_n307), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT38), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n295), .A2(new_n297), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n300), .A3(new_n282), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n306), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n298), .A2(new_n203), .A3(new_n300), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n524), .A2(new_n505), .A3(new_n512), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n198), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n512), .B1(new_n502), .B2(new_n505), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n541), .A2(new_n542), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n187), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n351), .A2(new_n659), .A3(new_n414), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n653), .A2(new_n624), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(KEYINPUT98), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n643), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n262), .ZN(G45));
  AOI211_X1 g479(.A(new_n659), .B(new_n624), .C1(new_n648), .C2(new_n649), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(new_n635), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n593), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(new_n593), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n491), .A2(new_n543), .A3(new_n666), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NAND3_X1  g487(.A1(new_n483), .A2(new_n198), .A3(new_n485), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(KEYINPUT100), .A3(new_n487), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n677), .A3(G469), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n580), .A3(new_n630), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n659), .B1(new_n648), .B2(new_n649), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n202), .A3(new_n593), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT101), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n418), .B1(new_n676), .B2(new_n678), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n595), .A2(new_n684), .A3(new_n685), .A4(new_n580), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND3_X1  g503(.A1(new_n606), .A2(new_n684), .A3(new_n580), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  INV_X1    g505(.A(new_n308), .ZN(new_n692));
  INV_X1    g506(.A(new_n415), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n543), .A2(new_n693), .A3(new_n625), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n684), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NOR2_X1   g510(.A1(new_n351), .A2(new_n414), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n512), .B1(new_n525), .B2(new_n534), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n531), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n533), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n699), .B1(new_n698), .B2(new_n531), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n538), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n579), .A3(new_n599), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n201), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n684), .A2(new_n681), .A3(new_n697), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND3_X1  g521(.A1(new_n625), .A2(new_n599), .A3(new_n703), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n684), .A2(new_n681), .A3(new_n671), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NOR2_X1   g525(.A1(new_n650), .A2(new_n659), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n477), .A2(G469), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n418), .B1(new_n713), .B2(new_n487), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n580), .A3(new_n671), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n187), .A2(new_n644), .A3(new_n714), .A4(new_n671), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n539), .A2(KEYINPUT103), .A3(new_n540), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n529), .A3(new_n542), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n539), .B2(new_n540), .ZN(new_n722));
  OAI211_X1 g536(.A(KEYINPUT42), .B(new_n579), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n718), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n644), .A2(new_n714), .A3(new_n671), .A4(new_n187), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n723), .A3(KEYINPUT104), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n717), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(KEYINPUT105), .B(new_n717), .C1(new_n725), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT106), .B(G131), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G33));
  NAND4_X1  g548(.A1(new_n712), .A2(new_n580), .A3(new_n636), .A4(new_n714), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(new_n469), .A2(new_n476), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n469), .A2(new_n476), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n487), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n741), .B2(new_n742), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n630), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n712), .B(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n590), .A2(new_n592), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n414), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n600), .A3(new_n625), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT44), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n641), .A2(new_n747), .A3(new_n748), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n426), .ZN(G39));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n745), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n487), .A3(new_n743), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n762), .B1(new_n764), .B2(new_n630), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n746), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(new_n762), .ZN(new_n767));
  INV_X1    g581(.A(new_n712), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n768), .A2(new_n543), .A3(new_n669), .A4(new_n670), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n767), .A2(new_n578), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n365), .ZN(G42));
  NOR3_X1   g585(.A1(new_n578), .A2(new_n418), .A3(new_n659), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n414), .A3(new_n749), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT110), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n679), .B(KEYINPUT49), .Z(new_n777));
  NOR4_X1   g591(.A1(new_n776), .A2(new_n777), .A3(new_n653), .A4(new_n658), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT111), .Z(new_n779));
  NAND3_X1  g593(.A1(new_n751), .A2(new_n752), .A3(new_n194), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n704), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n679), .A2(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n679), .A2(KEYINPUT114), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n418), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n748), .B(new_n781), .C1(new_n767), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n187), .B1(new_n645), .B2(new_n652), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n684), .A3(new_n781), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n194), .A2(new_n684), .A3(new_n712), .A4(new_n754), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n709), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n787), .A2(new_n684), .A3(new_n794), .A4(new_n781), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n684), .A2(new_n194), .A3(new_n712), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n658), .A2(new_n578), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n797), .A2(new_n413), .A3(new_n749), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n786), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n579), .B1(new_n721), .B2(new_n722), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n797), .A2(new_n802), .A3(new_n753), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT48), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n487), .A2(KEYINPUT100), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT79), .B1(new_n479), .B2(new_n463), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n484), .B1(new_n806), .B2(new_n482), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n486), .B1(new_n807), .B2(new_n198), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n678), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n681), .B(new_n630), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n781), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n797), .A2(new_n798), .ZN(new_n813));
  OAI221_X1 g627(.A(new_n190), .B1(new_n811), .B2(new_n812), .C1(new_n813), .C2(new_n594), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n801), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT116), .B1(new_n796), .B2(new_n799), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n709), .ZN(new_n818));
  INV_X1    g632(.A(new_n799), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n795), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n786), .A2(new_n817), .A3(KEYINPUT51), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n815), .B(new_n816), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n822), .B(KEYINPUT117), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n816), .B1(new_n828), .B2(new_n815), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n735), .B1(new_n708), .B2(new_n726), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n768), .A2(new_n632), .A3(new_n624), .A4(new_n635), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n693), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n732), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n683), .A2(new_n686), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n626), .A2(new_n602), .A3(new_n607), .A4(new_n581), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n706), .A2(new_n690), .A3(new_n695), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n671), .A2(new_n599), .A3(new_n625), .A4(new_n703), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n811), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT112), .B1(new_n840), .B2(new_n639), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n650), .A2(new_n660), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n615), .A2(new_n620), .A3(new_n635), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n658), .A3(new_n714), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n491), .A2(new_n543), .A3(new_n636), .A4(new_n666), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n710), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n841), .A2(new_n845), .A3(new_n848), .A4(new_n672), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n672), .A3(new_n710), .A4(new_n844), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n833), .A2(new_n834), .A3(new_n838), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n840), .A2(new_n639), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n844), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n852), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n732), .A2(new_n838), .A3(new_n857), .A4(new_n832), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(KEYINPUT54), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n834), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n706), .A2(new_n690), .A3(new_n695), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n728), .A2(new_n687), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n728), .A2(new_n862), .A3(new_n687), .A4(KEYINPUT113), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n626), .A2(new_n581), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n602), .A4(new_n607), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n852), .B2(new_n849), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n832), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n860), .B1(KEYINPUT54), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n827), .A2(new_n829), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n779), .B1(new_n874), .B2(new_n875), .ZN(G75));
  XOR2_X1   g690(.A(new_n296), .B(KEYINPUT55), .Z(new_n877));
  XOR2_X1   g691(.A(new_n295), .B(KEYINPUT119), .Z(new_n878));
  AOI21_X1  g692(.A(new_n198), .B1(new_n861), .B2(new_n871), .ZN(new_n879));
  AOI211_X1 g693(.A(KEYINPUT56), .B(new_n878), .C1(new_n879), .C2(G210), .ZN(new_n880));
  INV_X1    g694(.A(new_n878), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n199), .A2(G952), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT120), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(G210), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n889), .B(new_n198), .C1(new_n861), .C2(new_n871), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n878), .B1(new_n890), .B2(KEYINPUT56), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n883), .A3(new_n881), .ZN(new_n892));
  INV_X1    g706(.A(new_n877), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n885), .A2(new_n888), .A3(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n742), .A2(KEYINPUT57), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n742), .A2(KEYINPUT57), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n807), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n741), .B(KEYINPUT121), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n879), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n886), .B1(new_n901), .B2(new_n903), .ZN(G54));
  NAND3_X1  g718(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n905));
  INV_X1    g719(.A(new_n404), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n886), .ZN(G60));
  AND2_X1   g723(.A1(new_n585), .A2(new_n589), .ZN(new_n910));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n912), .C1(new_n898), .C2(new_n899), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n873), .B2(new_n912), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n887), .A3(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT122), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n872), .A2(new_n618), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n872), .A2(new_n919), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n888), .B(new_n920), .C1(new_n921), .C2(new_n569), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n920), .B2(KEYINPUT123), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G66));
  AOI21_X1  g738(.A(new_n199), .B1(new_n196), .B2(G224), .ZN(new_n925));
  INV_X1    g739(.A(new_n838), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n199), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n881), .B1(G898), .B2(new_n199), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  NAND2_X1  g744(.A1(G227), .A2(G900), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n633), .A2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT126), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n770), .A2(new_n757), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n841), .A2(new_n848), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n672), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n747), .A2(new_n641), .A3(new_n842), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n732), .B(new_n735), .C1(new_n939), .C2(new_n802), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n941), .B2(G953), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n497), .A2(new_n501), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n393), .A2(new_n394), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n664), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(KEYINPUT62), .A3(new_n672), .A4(new_n937), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n938), .B2(new_n664), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n642), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n605), .A2(new_n594), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n580), .A3(new_n712), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n935), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n951), .A2(new_n957), .A3(new_n935), .A4(new_n954), .ZN(new_n958));
  AOI21_X1  g772(.A(G953), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n932), .B(new_n946), .C1(new_n959), .C2(new_n945), .ZN(new_n960));
  INV_X1    g774(.A(new_n945), .ZN(new_n961));
  OAI211_X1 g775(.A(G953), .B(new_n931), .C1(new_n942), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(G72));
  NOR2_X1   g777(.A1(new_n506), .A2(new_n511), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n936), .A2(new_n926), .A3(new_n940), .A4(new_n938), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n513), .ZN(new_n970));
  INV_X1    g784(.A(new_n530), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT127), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n968), .B(new_n972), .C1(KEYINPUT127), .C2(new_n970), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n854), .A2(new_n859), .A3(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n969), .B(new_n974), .C1(G952), .C2(new_n199), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n956), .A2(new_n838), .A3(new_n958), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n967), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n656), .B2(new_n977), .ZN(G57));
endmodule


