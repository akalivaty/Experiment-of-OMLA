//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n668, new_n671, new_n673, new_n674, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT65), .Z(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n463));
  NAND4_X1  g038(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g052(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G112), .B2(new_n467), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n460), .A2(new_n463), .A3(new_n462), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n482), .A2(new_n486), .A3(new_n467), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n482), .B2(new_n467), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n489), .B2(G136), .ZN(G162));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n460), .A2(new_n462), .A3(new_n497), .A4(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT3), .B(G2104), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n497), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n499), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n513), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI211_X1 g090(.A(new_n507), .B(new_n515), .C1(new_n510), .C2(new_n512), .ZN(new_n516));
  OAI21_X1  g091(.A(G62), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(G88), .B(new_n524), .C1(new_n514), .C2(new_n516), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n515), .B1(new_n527), .B2(new_n520), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n505), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT72), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n534), .B2(new_n515), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT72), .B(G543), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n532), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n518), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n529), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n523), .B1(new_n535), .B2(new_n538), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(G88), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT73), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n531), .A2(new_n545), .ZN(G166));
  NAND2_X1  g121(.A1(new_n543), .A2(G89), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n535), .A2(new_n538), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n548), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n552));
  AOI22_X1  g127(.A1(G51), .A2(new_n528), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n547), .A2(new_n549), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  AND2_X1   g130(.A1(new_n548), .A2(G64), .ZN(new_n556));
  AND2_X1   g131(.A1(G77), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT74), .B(G90), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI211_X1 g135(.A(new_n523), .B(new_n560), .C1(new_n535), .C2(new_n538), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n528), .A2(G52), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n548), .A2(new_n524), .A3(new_n559), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n566), .B2(new_n563), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n558), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(new_n573), .A3(new_n558), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(G171));
  AOI22_X1  g150(.A1(new_n543), .A2(G81), .B1(G43), .B2(new_n528), .ZN(new_n576));
  INV_X1    g151(.A(G56), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n535), .B2(new_n538), .ZN(new_n578));
  NAND2_X1  g153(.A1(G68), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n576), .B2(new_n581), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G860), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g163(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g164(.A1(G1), .A2(G3), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT8), .ZN(new_n591));
  NAND4_X1  g166(.A1(G319), .A2(G483), .A3(G661), .A4(new_n591), .ZN(G188));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  INV_X1    g168(.A(G65), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n535), .B2(new_n538), .ZN(new_n595));
  AND2_X1   g170(.A1(G78), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n543), .A2(G91), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT9), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n528), .B2(G53), .ZN(new_n602));
  OAI211_X1 g177(.A(G53), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(KEYINPUT9), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n528), .A2(new_n601), .A3(G53), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(KEYINPUT9), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT79), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n593), .B1(new_n599), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(new_n597), .A3(new_n598), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n612), .ZN(G299));
  INV_X1    g188(.A(G171), .ZN(G301));
  AND3_X1   g189(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT73), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT73), .B1(new_n541), .B2(new_n544), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT81), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n531), .A2(new_n545), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n617), .A2(new_n619), .ZN(G303));
  NOR2_X1   g195(.A1(new_n514), .A2(new_n516), .ZN(new_n621));
  INV_X1    g196(.A(G74), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G49), .B2(new_n528), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n543), .A2(G87), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n625), .A2(KEYINPUT82), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(KEYINPUT82), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(G288));
  OAI211_X1 g203(.A(G86), .B(new_n524), .C1(new_n514), .C2(new_n516), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n528), .A2(G48), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n632));
  INV_X1    g207(.A(G61), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n535), .B2(new_n538), .ZN(new_n634));
  AND2_X1   g209(.A1(G73), .A2(G543), .ZN(new_n635));
  OAI21_X1  g210(.A(G651), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n631), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(KEYINPUT83), .B(G651), .C1(new_n634), .C2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(G305));
  AOI22_X1  g214(.A1(new_n548), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(new_n506), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(G47), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n543), .A2(G85), .B1(new_n528), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(G290));
  INV_X1    g219(.A(G868), .ZN(new_n645));
  NOR2_X1   g220(.A1(G301), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n548), .A2(G92), .A3(new_n524), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n543), .A2(KEYINPUT10), .A3(G92), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n528), .A2(G54), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n548), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n506), .ZN(new_n654));
  OAI21_X1  g229(.A(KEYINPUT85), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(G79), .A2(G543), .ZN(new_n656));
  INV_X1    g231(.A(G66), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n621), .B2(new_n657), .ZN(new_n658));
  AOI22_X1  g233(.A1(new_n658), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n649), .A2(new_n650), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n646), .B1(new_n665), .B2(new_n645), .ZN(G284));
  AOI21_X1  g241(.A(new_n646), .B1(new_n665), .B2(new_n645), .ZN(G321));
  NAND2_X1  g242(.A1(G299), .A2(new_n645), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n645), .B2(G168), .ZN(G297));
  OAI21_X1  g244(.A(new_n668), .B1(new_n645), .B2(G168), .ZN(G280));
  INV_X1    g245(.A(G559), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n665), .B1(new_n671), .B2(G860), .ZN(G148));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G868), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G868), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g250(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g251(.A(new_n483), .ZN(new_n677));
  OAI21_X1  g252(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G111), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n678), .A2(new_n679), .B1(new_n681), .B2(G2105), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n677), .A2(G123), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n489), .B2(G135), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(G2096), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(G2096), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT12), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT13), .ZN(new_n691));
  NAND2_X1  g266(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n691), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(KEYINPUT87), .B2(G2100), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n693), .B1(new_n695), .B2(new_n692), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n687), .A2(new_n688), .A3(new_n696), .ZN(G156));
  XNOR2_X1  g272(.A(G2427), .B(G2438), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2430), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT15), .B(G2435), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(KEYINPUT14), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  XOR2_X1   g279(.A(G1341), .B(G1348), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G2451), .B(G2454), .Z(new_n707));
  XNOR2_X1  g282(.A(G2443), .B(G2446), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n706), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n713), .A3(G14), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G401));
  INV_X1    g290(.A(KEYINPUT18), .ZN(new_n716));
  XOR2_X1   g291(.A(G2084), .B(G2090), .Z(new_n717));
  XNOR2_X1  g292(.A(G2067), .B(G2678), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT17), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2100), .ZN(new_n723));
  XOR2_X1   g298(.A(G2072), .B(G2078), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n719), .B2(KEYINPUT18), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2096), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n723), .B(new_n726), .ZN(G227));
  XOR2_X1   g302(.A(G1971), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT19), .ZN(new_n729));
  XOR2_X1   g304(.A(G1956), .B(G2474), .Z(new_n730));
  XOR2_X1   g305(.A(G1961), .B(G1966), .Z(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT20), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n730), .A2(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n729), .A2(new_n732), .A3(new_n735), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(G1991), .B(G1996), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(G1981), .B(G1986), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n745), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(G229));
  MUX2_X1   g323(.A(G23), .B(G288), .S(G16), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT33), .B(G1976), .Z(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G6), .B(G305), .S(G16), .Z(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT32), .B(G1981), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G22), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G166), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1971), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n750), .B2(new_n752), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT34), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n757), .A2(new_n765), .A3(new_n762), .ZN(new_n766));
  INV_X1    g341(.A(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G25), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n489), .A2(G131), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G107), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n677), .B2(G119), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n768), .B1(new_n775), .B2(new_n767), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT35), .B(G1991), .Z(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n776), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT94), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n758), .A2(G24), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  INV_X1    g358(.A(G290), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n758), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n781), .B1(new_n785), .B2(G1986), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G1986), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n764), .A2(new_n766), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n789), .A2(KEYINPUT94), .A3(new_n780), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n780), .A2(KEYINPUT94), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n764), .A2(new_n791), .A3(new_n766), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT104), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G34), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n767), .B1(new_n795), .B2(G34), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n474), .A2(new_n767), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2084), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n767), .A2(G32), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n489), .A2(G141), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  NAND3_X1  g379(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n677), .B2(G129), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n800), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n767), .A2(G33), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n489), .A2(G139), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n500), .A2(G127), .ZN(new_n814));
  INV_X1    g389(.A(G115), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n459), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n817));
  NAND2_X1  g392(.A1(G103), .A2(G2104), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n816), .A2(G2105), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n812), .B1(new_n822), .B2(new_n767), .ZN(new_n823));
  INV_X1    g398(.A(G2072), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n811), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT101), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n758), .A2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G168), .B2(new_n758), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT102), .Z(new_n831));
  INV_X1    g406(.A(G1966), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT103), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n809), .A2(new_n810), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n686), .A2(new_n767), .ZN(new_n837));
  NOR2_X1   g412(.A1(G27), .A2(G29), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G164), .B2(G29), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(G2078), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(G2078), .ZN(new_n841));
  INV_X1    g416(.A(G28), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT30), .ZN(new_n843));
  AOI21_X1  g418(.A(G29), .B1(new_n842), .B2(KEYINPUT30), .ZN(new_n844));
  OR2_X1    g419(.A1(KEYINPUT31), .A2(G11), .ZN(new_n845));
  NAND2_X1  g420(.A1(KEYINPUT31), .A2(G11), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n798), .A2(new_n799), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n840), .A2(new_n841), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NOR4_X1   g424(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n758), .A2(G5), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G171), .B2(new_n758), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(G1961), .Z(new_n853));
  NAND3_X1  g428(.A1(new_n834), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n794), .B1(new_n828), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n827), .B(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n834), .A2(new_n850), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(KEYINPUT104), .A3(new_n858), .A4(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n758), .A2(G4), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n665), .B2(new_n758), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT96), .B(G1348), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT95), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n767), .A2(G26), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT28), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n489), .A2(new_n867), .A3(G140), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n487), .A2(new_n488), .ZN(new_n869));
  INV_X1    g444(.A(G140), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n873));
  OR3_X1    g448(.A1(KEYINPUT99), .A2(G104), .A3(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT99), .B1(G104), .B2(G2105), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n677), .B2(G128), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n866), .B1(new_n878), .B2(new_n767), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT100), .B(G2067), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(G16), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n758), .A2(G20), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT23), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(G1956), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n758), .A2(G19), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT97), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n576), .A2(new_n581), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT77), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n583), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n892), .B2(G16), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(G1341), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n767), .A2(G35), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(G162), .B2(new_n767), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT29), .B(G2090), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n887), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n864), .A2(new_n881), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n855), .A2(new_n859), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n793), .A2(new_n901), .ZN(G311));
  AND2_X1   g477(.A1(new_n859), .A2(new_n900), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(new_n855), .A3(new_n790), .A4(new_n792), .ZN(G150));
  AOI22_X1  g479(.A1(new_n548), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(new_n506), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n543), .A2(G93), .B1(G55), .B2(new_n528), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT106), .B(G860), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n892), .A2(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n890), .B2(new_n908), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n665), .A2(G559), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n915), .B(new_n916), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT39), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n918), .B2(new_n909), .ZN(G145));
  INV_X1    g494(.A(new_n808), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n822), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n813), .A2(new_n821), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n808), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n925));
  INV_X1    g500(.A(G118), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(G2105), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n677), .B2(G130), .ZN(new_n928));
  INV_X1    g503(.A(G142), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n869), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(new_n690), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n923), .A3(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n878), .A2(G164), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n872), .A2(new_n877), .ZN(new_n937));
  INV_X1    g512(.A(G164), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n774), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n774), .B1(new_n936), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n939), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n937), .A2(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n775), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n940), .A3(new_n934), .A4(new_n932), .ZN(new_n947));
  XNOR2_X1  g522(.A(G162), .B(new_n474), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(new_n685), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n943), .B2(new_n947), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT40), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(G395));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n659), .A2(new_n660), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n610), .A2(new_n612), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n599), .A2(new_n593), .A3(new_n609), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(new_n660), .B2(new_n659), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n957), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n610), .B2(new_n612), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n660), .A4(new_n659), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n914), .B1(new_n665), .B2(new_n671), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n665), .A2(new_n671), .A3(new_n914), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n972), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n965), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(new_n970), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT42), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(G305), .B(G288), .ZN(new_n978));
  XNOR2_X1  g553(.A(G166), .B(G290), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n968), .B(new_n963), .C1(new_n974), .C2(new_n970), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n971), .A2(new_n972), .A3(new_n965), .A4(new_n964), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n977), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n977), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g564(.A(G868), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n908), .A2(new_n645), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(G295));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n991), .ZN(G331));
  AND2_X1   g568(.A1(new_n576), .A2(new_n581), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n994), .A2(new_n906), .A3(new_n907), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n892), .B2(new_n908), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n573), .B1(new_n572), .B2(new_n558), .ZN(new_n998));
  OAI21_X1  g573(.A(G168), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n569), .A2(G286), .A3(new_n574), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n969), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n914), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n975), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n982), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n951), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT109), .B(new_n966), .C1(new_n959), .C2(new_n962), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n964), .A2(KEYINPUT41), .A3(new_n965), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT109), .B1(new_n975), .B2(new_n966), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n1012), .A2(new_n1013), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n982), .B1(new_n1014), .B2(new_n1007), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n983), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n951), .A4(new_n1008), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(KEYINPUT44), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT110), .A4(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1009), .B1(new_n1017), .B2(new_n983), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n1019), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1009), .A2(new_n1015), .A3(KEYINPUT43), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(G397));
  OR2_X1    g606(.A1(G288), .A2(G1976), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n500), .A2(new_n1035), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1036), .B2(new_n495), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n468), .A2(G40), .A3(new_n473), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n637), .B2(new_n638), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n636), .A2(new_n632), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n629), .A2(new_n630), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1042), .A3(new_n638), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n637), .A2(KEYINPUT117), .A3(new_n1042), .A4(new_n638), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1041), .B1(new_n1050), .B2(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1052), .B(new_n1043), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1033), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT119), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1041), .B(KEYINPUT118), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1041), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1043), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1061), .B2(new_n1052), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n624), .B(G1976), .C1(new_n626), .C2(new_n627), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(KEYINPUT116), .A3(new_n1041), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G288), .A2(new_n1064), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1041), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1041), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1062), .A2(new_n1063), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n617), .A2(G8), .A3(new_n619), .ZN(new_n1076));
  AND2_X1   g651(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  AOI21_X1  g655(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n1081));
  INV_X1    g656(.A(G40), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n472), .ZN(new_n1083));
  NOR2_X1   g658(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1036), .B2(new_n495), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT45), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(G164), .B2(G1384), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT45), .B(new_n1034), .C1(new_n1036), .C2(new_n495), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT113), .B(G1971), .ZN(new_n1091));
  AOI22_X1  g666(.A1(KEYINPUT114), .A2(new_n1086), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1040), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1077), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n617), .A2(G8), .A3(new_n619), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1078), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1057), .A2(new_n1058), .B1(new_n1075), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1086), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1040), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(KEYINPUT120), .A3(new_n1086), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1078), .A2(new_n1097), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1079), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1038), .B1(new_n1037), .B2(new_n1087), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1089), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n606), .B2(new_n607), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n599), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n611), .A2(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1110), .A2(new_n1113), .A3(new_n1117), .A4(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n659), .A2(new_n661), .A3(new_n660), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G2067), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1108), .A2(new_n862), .B1(new_n1039), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n655), .A2(new_n1127), .A3(new_n662), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n583), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(G1996), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n499), .A2(new_n503), .ZN(new_n1132));
  INV_X1    g707(.A(new_n495), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1384), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1134), .B2(KEYINPUT45), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1083), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  AOI22_X1  g712(.A1(new_n1111), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT59), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1083), .B1(new_n1134), .B2(KEYINPUT45), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1131), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1089), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n586), .A2(new_n1144), .A3(KEYINPUT123), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1126), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n663), .A3(KEYINPUT60), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1121), .A2(new_n1129), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1119), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1126), .B1(new_n655), .B2(new_n662), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1120), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G2078), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1111), .A2(new_n1155), .A3(new_n1089), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT124), .B(G1961), .Z(new_n1158));
  AOI22_X1  g733(.A1(new_n1156), .A2(new_n1157), .B1(new_n1108), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1141), .A2(new_n1160), .B1(KEYINPUT45), .B2(new_n1134), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1111), .A2(KEYINPUT121), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1157), .A2(G2078), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n569), .A2(KEYINPUT54), .A3(new_n574), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT54), .B1(new_n569), .B2(new_n574), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n997), .B2(new_n998), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n569), .A2(KEYINPUT54), .A3(new_n574), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1089), .A3(new_n1173), .A4(new_n1163), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1170), .A2(new_n1171), .A3(new_n1159), .A4(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1120), .A2(KEYINPUT61), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1168), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1107), .A2(new_n1154), .A3(new_n1177), .A4(new_n1075), .ZN(new_n1178));
  AOI21_X1  g753(.A(G1966), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1108), .A2(G2084), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g756(.A(KEYINPUT51), .B(new_n1040), .C1(new_n1181), .C2(G168), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1040), .B1(new_n1181), .B2(G168), .ZN(new_n1183));
  OAI21_X1  g758(.A(G286), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1185), .B2(KEYINPUT51), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1100), .B1(new_n1178), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1078), .A2(new_n1097), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g765(.A(G8), .B(G168), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1075), .A2(new_n1098), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1098), .A2(KEYINPUT63), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1094), .B1(new_n1078), .B2(new_n1097), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1195), .A2(new_n1191), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1193), .A2(new_n1194), .B1(new_n1197), .B2(new_n1075), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT126), .B1(new_n1187), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1061), .A2(new_n1052), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n1063), .A3(new_n1041), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1074), .A2(new_n1067), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1201), .A2(new_n1190), .A3(new_n1202), .A4(new_n1098), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1194), .B1(new_n1203), .B2(new_n1191), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1197), .A2(new_n1075), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1185), .A2(KEYINPUT51), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1182), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1203), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1168), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1212), .B1(new_n1153), .B2(new_n1150), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1206), .A2(new_n1207), .A3(new_n1214), .A4(new_n1100), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1210), .A2(KEYINPUT62), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1186), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(G301), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1216), .A2(new_n1211), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1199), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n937), .B(new_n1125), .ZN(new_n1222));
  INV_X1    g797(.A(G1996), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1223), .B2(new_n920), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1088), .A2(new_n1038), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1223), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT112), .ZN(new_n1227));
  AOI22_X1  g802(.A1(new_n1224), .A2(new_n1225), .B1(new_n920), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n775), .A2(new_n777), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n774), .A2(new_n778), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1225), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1225), .ZN(new_n1233));
  NOR2_X1   g808(.A1(G290), .A2(G1986), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT111), .ZN(new_n1235));
  NAND2_X1  g810(.A1(G290), .A2(G1986), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1221), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1235), .A2(new_n1233), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1240), .B(KEYINPUT48), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1233), .B1(new_n1222), .B2(new_n920), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1227), .B1(KEYINPUT127), .B2(KEYINPUT46), .ZN(new_n1243));
  NAND2_X1  g818(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1244));
  MUX2_X1   g819(.A(new_n1227), .B(new_n1243), .S(new_n1244), .Z(new_n1245));
  NOR2_X1   g820(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT47), .ZN(new_n1247));
  NOR2_X1   g822(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1242), .A2(new_n1245), .A3(KEYINPUT47), .ZN(new_n1249));
  OAI22_X1  g824(.A1(new_n1232), .A2(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n878), .A2(new_n1125), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1233), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g828(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1239), .A2(new_n1254), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1257));
  INV_X1    g831(.A(G319), .ZN(new_n1258));
  OR2_X1    g832(.A1(G227), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g833(.A(new_n1259), .B1(new_n746), .B2(new_n747), .ZN(new_n1260));
  OAI211_X1 g834(.A(new_n1260), .B(new_n714), .C1(new_n952), .C2(new_n953), .ZN(new_n1261));
  NOR2_X1   g835(.A1(new_n1257), .A2(new_n1261), .ZN(G308));
  AND2_X1   g836(.A1(new_n1260), .A2(new_n714), .ZN(new_n1263));
  OAI221_X1 g837(.A(new_n1263), .B1(new_n952), .B2(new_n953), .C1(new_n1028), .C2(new_n1029), .ZN(G225));
endmodule


