//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n209), .B2(new_n211), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n206), .B(new_n207), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT81), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n210), .A2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n208), .A2(G141gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT79), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n206), .A4(new_n207), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT2), .B1(new_n209), .B2(new_n211), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT78), .B1(new_n225), .B2(new_n207), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n205), .A2(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231));
  XNOR2_X1  g030(.A(G141gat), .B(G148gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239));
  INV_X1    g038(.A(G120gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(G113gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(G120gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n241), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n237), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n234), .B1(new_n216), .B2(new_n223), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n252), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n254), .B2(new_n255), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT3), .B(new_n234), .C1(new_n216), .C2(new_n223), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n252), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n253), .A2(new_n202), .ZN(new_n265));
  OAI211_X1 g064(.A(KEYINPUT5), .B(new_n257), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n203), .A2(KEYINPUT5), .ZN(new_n267));
  OAI221_X1 g066(.A(new_n267), .B1(new_n263), .B2(new_n261), .C1(new_n258), .C2(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT0), .B(G57gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G85gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G1gat), .B(G29gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n273), .A3(new_n268), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT86), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n273), .B1(new_n266), .B2(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT6), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n275), .A2(new_n282), .A3(new_n276), .A4(new_n277), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT27), .B(G183gat), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT66), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT65), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  OR3_X1    g092(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n295), .A2(KEYINPUT67), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT67), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n296), .A2(KEYINPUT24), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n287), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT24), .A3(new_n296), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n306), .A4(new_n292), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n292), .A2(new_n306), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n310), .A2(new_n302), .A3(KEYINPUT25), .A4(new_n303), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n299), .B2(new_n312), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n314), .B(KEYINPUT75), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G211gat), .A2(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT73), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n326), .A3(new_n322), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(new_n329), .A3(new_n325), .A4(new_n327), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT74), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n319), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n332), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n338), .B(new_n339), .C1(new_n317), .C2(new_n315), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  INV_X1    g140(.A(G64gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G92gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n317), .A2(new_n315), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n313), .B2(new_n319), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n349), .A2(new_n339), .B1(new_n336), .B2(new_n320), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT37), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n337), .A2(new_n340), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT37), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT38), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n351), .A2(new_n355), .A3(new_n356), .A4(new_n345), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n284), .A2(new_n285), .A3(new_n347), .A4(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n278), .A2(KEYINPUT86), .B1(KEYINPUT6), .B2(new_n280), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(new_n347), .A3(new_n283), .A4(new_n357), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT87), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n345), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n353), .A2(new_n354), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT38), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n262), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n236), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G228gat), .ZN(new_n372));
  INV_X1    g171(.A(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n254), .B2(new_n262), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n371), .B(new_n374), .C1(new_n375), .C2(new_n335), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n339), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n379), .B2(new_n371), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n367), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT31), .ZN(new_n383));
  INV_X1    g182(.A(G50gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n374), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n224), .A2(new_n262), .A3(new_n235), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n339), .B1(new_n388), .B2(new_n368), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n254), .B1(new_n262), .B2(new_n369), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(G22gat), .A3(new_n376), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n381), .A2(new_n386), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT82), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n381), .A2(new_n392), .A3(new_n395), .A4(new_n386), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n367), .A2(KEYINPUT83), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n391), .A2(new_n376), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n391), .B2(new_n376), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n385), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT84), .ZN(new_n402));
  INV_X1    g201(.A(new_n398), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n377), .B2(new_n380), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n391), .A2(new_n376), .A3(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n385), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n397), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n406), .B2(new_n385), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT84), .B(new_n386), .C1(new_n404), .C2(new_n405), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n396), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n346), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n352), .A2(new_n345), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n347), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n264), .A2(new_n203), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n253), .A2(new_n256), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(KEYINPUT39), .C1(new_n203), .C2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n273), .C1(KEYINPUT39), .C2(new_n428), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n280), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n366), .A2(new_n418), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT70), .B1(new_n249), .B2(new_n251), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n252), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n288), .B(KEYINPUT28), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n295), .A2(KEYINPUT67), .A3(new_n296), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n295), .A2(new_n296), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n309), .A2(new_n311), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n442), .B(new_n445), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G227gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(new_n373), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n299), .A2(new_n443), .A3(new_n252), .A4(new_n312), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT71), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n453), .A2(KEYINPUT71), .A3(new_n455), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n440), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n455), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n441), .B(new_n444), .C1(new_n299), .C2(new_n312), .ZN(new_n466));
  INV_X1    g265(.A(new_n456), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT34), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n459), .B2(new_n460), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n469), .A3(new_n471), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n474), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n463), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT72), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n421), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n491), .A2(new_n492), .B1(new_n424), .B2(new_n425), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n278), .A2(new_n281), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n494), .C1(new_n492), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n417), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n436), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n410), .B1(new_n397), .B2(new_n409), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n415), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n482), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT35), .B1(new_n503), .B2(new_n495), .ZN(new_n504));
  AOI211_X1 g303(.A(KEYINPUT35), .B(new_n482), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n284), .A2(new_n427), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT88), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n483), .C1(new_n411), .C2(new_n416), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n359), .A2(new_n283), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n426), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n504), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(KEYINPUT15), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  AND2_X1   g331(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(KEYINPUT17), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n521), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n532), .B(new_n521), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n536), .B(KEYINPUT13), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G113gat), .B(G141gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT98), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G120gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n208), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n559), .B(KEYINPUT94), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n567), .B2(new_n344), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n562), .A2(new_n565), .A3(new_n572), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n573), .ZN(new_n574));
  OR3_X1    g373(.A1(new_n569), .A2(KEYINPUT95), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n342), .A2(G57gat), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT90), .B(G57gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n579), .B2(new_n342), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n573), .A3(new_n571), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n596), .B(new_n590), .C1(new_n576), .C2(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n576), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT99), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n596), .B1(new_n576), .B2(new_n595), .ZN(new_n603));
  INV_X1    g402(.A(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n558), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n605), .A3(new_n557), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n553), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n521), .B1(new_n589), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT92), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n589), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n617), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n622), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n534), .A2(new_n575), .A3(new_n574), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n576), .A2(new_n532), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT93), .Z(new_n631));
  OAI211_X1 g430(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G190gat), .B(G218gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n629), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640));
  INV_X1    g439(.A(new_n633), .ZN(new_n641));
  OR3_X1    g440(.A1(new_n632), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n634), .A2(new_n640), .A3(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n612), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n515), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n494), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n427), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n517), .A2(new_n520), .ZN(new_n653));
  NOR2_X1   g452(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n655));
  NOR4_X1   g454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(G8gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n648), .B2(new_n483), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n490), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(G15gat), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n647), .A2(new_n418), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT102), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n666), .B(new_n668), .ZN(G1327gat));
  AOI21_X1  g468(.A(new_n644), .B1(new_n499), .B2(new_n514), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n612), .A2(new_n626), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n524), .A3(new_n649), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n510), .B1(new_n509), .B2(new_n512), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n506), .A2(KEYINPUT88), .A3(new_n502), .A4(new_n508), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n677), .A2(new_n678), .A3(new_n504), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n677), .B2(new_n504), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n499), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n644), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT44), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n684), .B(new_n644), .C1(new_n499), .C2(new_n514), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n671), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n494), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n674), .B1(new_n689), .B2(new_n524), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n525), .A3(new_n427), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT46), .Z(new_n692));
  NOR3_X1   g491(.A1(new_n687), .A2(new_n426), .A3(new_n688), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n525), .B2(new_n693), .ZN(G1329gat));
  NOR4_X1   g493(.A1(new_n683), .A2(new_n685), .A3(new_n490), .A4(new_n688), .ZN(new_n695));
  INV_X1    g494(.A(G43gat), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n696), .A3(new_n483), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI221_X1 g500(.A(new_n698), .B1(KEYINPUT104), .B2(KEYINPUT47), .C1(new_n695), .C2(new_n696), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  INV_X1    g502(.A(new_n435), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n362), .B2(new_n365), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n497), .B1(new_n705), .B2(new_n418), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n514), .A2(KEYINPUT103), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n677), .A2(new_n678), .A3(new_n504), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n684), .B1(new_n709), .B2(new_n644), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n670), .A2(KEYINPUT44), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n417), .A3(new_n671), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT105), .B1(new_n712), .B2(G50gat), .ZN(new_n713));
  AND4_X1   g512(.A1(new_n384), .A2(new_n670), .A3(new_n417), .A4(new_n671), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n712), .B2(G50gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI221_X4 g516(.A(new_n714), .B1(KEYINPUT105), .B2(KEYINPUT48), .C1(new_n712), .C2(G50gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n610), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n550), .A2(new_n552), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n645), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n709), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n494), .B(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n579), .ZN(G1332gat));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n426), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  INV_X1    g532(.A(G71gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n728), .B2(new_n482), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n681), .A2(G71gat), .A3(new_n610), .A4(new_n722), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n490), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(KEYINPUT107), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n736), .A2(new_n739), .A3(new_n490), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n735), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT50), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n735), .B(new_n743), .C1(new_n738), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n417), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n626), .A2(new_n721), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n681), .A2(new_n682), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n751), .A2(new_n567), .A3(new_n649), .A4(new_n610), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n710), .A2(new_n610), .A3(new_n711), .A4(new_n748), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n494), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1336gat));
  NOR3_X1   g554(.A1(new_n426), .A2(G92gat), .A3(new_n720), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G92gat), .B1(new_n753), .B2(new_n426), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n749), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n749), .B2(KEYINPUT109), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n756), .B(KEYINPUT108), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n686), .A2(new_n427), .A3(new_n610), .A4(new_n748), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(G1337gat));
  NOR2_X1   g567(.A1(new_n482), .A2(G99gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n610), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G99gat), .B1(new_n753), .B2(new_n490), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1338gat));
  NOR3_X1   g571(.A1(new_n418), .A2(G106gat), .A3(new_n720), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT111), .Z(new_n774));
  AOI21_X1  g573(.A(KEYINPUT53), .B1(new_n751), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n686), .A2(new_n417), .A3(new_n610), .A4(new_n748), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n774), .B(KEYINPUT112), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n763), .A2(new_n779), .B1(new_n776), .B2(G106gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(new_n626), .ZN(new_n783));
  INV_X1    g582(.A(new_n609), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n608), .B(KEYINPUT54), .C1(new_n601), .C2(new_n599), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n599), .A2(new_n786), .A3(new_n601), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n558), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n787), .B2(new_n558), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT55), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n792), .B(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n784), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n721), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n539), .A2(new_n540), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT114), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n535), .A2(new_n536), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n548), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n552), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n610), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n682), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n682), .A2(new_n794), .A3(new_n800), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n783), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n722), .A2(new_n720), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(new_n426), .A3(new_n725), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n502), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n243), .A3(new_n721), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n427), .A2(new_n494), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n502), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n553), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(G1340gat));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n240), .A3(new_n610), .ZN(new_n814));
  OAI21_X1  g613(.A(G120gat), .B1(new_n811), .B2(new_n720), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT115), .Z(G1341gat));
  INV_X1    g616(.A(G127gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n811), .A2(new_n818), .A3(new_n783), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n808), .A2(new_n626), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n818), .ZN(G1342gat));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n808), .A2(new_n822), .A3(new_n682), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT56), .Z(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n811), .B2(new_n644), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1343gat));
  NOR2_X1   g625(.A1(new_n489), .A2(new_n418), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n807), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(new_n210), .A3(new_n721), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n791), .A2(new_n793), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT116), .A3(new_n609), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n721), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n801), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n803), .B1(new_n836), .B2(new_n644), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n805), .B1(new_n837), .B2(new_n626), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n831), .B1(new_n838), .B2(new_n417), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n831), .A3(new_n417), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n490), .A2(new_n810), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n839), .A2(new_n843), .A3(new_n553), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n830), .B1(new_n210), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n839), .A2(new_n843), .A3(KEYINPUT117), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  INV_X1    g646(.A(new_n805), .ZN(new_n848));
  INV_X1    g647(.A(new_n803), .ZN(new_n849));
  INV_X1    g648(.A(new_n801), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n553), .B1(new_n794), .B2(KEYINPUT116), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n853), .B2(new_n682), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n848), .B1(new_n854), .B2(new_n783), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n418), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n418), .B1(new_n804), .B2(new_n805), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n841), .B1(new_n857), .B2(new_n831), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n847), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n721), .B1(new_n846), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n829), .B1(new_n860), .B2(G141gat), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n845), .B1(new_n861), .B2(new_n862), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n828), .A2(new_n208), .A3(new_n610), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n857), .A2(new_n831), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n854), .A2(new_n783), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n418), .B1(new_n867), .B2(new_n805), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(new_n831), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n841), .B(KEYINPUT118), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n610), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n208), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n869), .A2(KEYINPUT119), .A3(new_n610), .A4(new_n870), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT117), .B1(new_n839), .B2(new_n843), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n856), .A2(new_n847), .A3(new_n858), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n720), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(KEYINPUT59), .A3(new_n208), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n864), .B1(new_n875), .B2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n828), .B2(new_n626), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n783), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(G155gat), .ZN(G1346gat));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n682), .B1(new_n846), .B2(new_n859), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT80), .B(G162gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n828), .A2(new_n888), .A3(new_n682), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n644), .B1(new_n876), .B2(new_n877), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n884), .B(new_n889), .C1(new_n891), .C2(new_n888), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n890), .A2(new_n893), .ZN(G1347gat));
  AOI21_X1  g693(.A(new_n649), .B1(new_n804), .B2(new_n805), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(new_n502), .A3(new_n427), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT121), .Z(new_n897));
  INV_X1    g696(.A(G169gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n898), .A3(new_n721), .ZN(new_n899));
  INV_X1    g698(.A(new_n806), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n725), .A2(new_n426), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n503), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n553), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n897), .B2(new_n610), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n720), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(G176gat), .B2(new_n907), .ZN(G1349gat));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  OAI21_X1  g709(.A(G183gat), .B1(new_n903), .B2(new_n783), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n286), .A3(new_n626), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n910), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1350gat));
  AOI21_X1  g717(.A(new_n287), .B1(new_n902), .B2(new_n682), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT61), .Z(new_n920));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n287), .A3(new_n682), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  AND3_X1   g721(.A1(new_n895), .A2(new_n427), .A3(new_n827), .ZN(new_n923));
  INV_X1    g722(.A(G197gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n721), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n901), .A2(new_n489), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT124), .Z(new_n927));
  AND3_X1   g726(.A1(new_n869), .A2(new_n721), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n924), .ZN(G1352gat));
  INV_X1    g728(.A(G204gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n930), .A3(new_n610), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  AND3_X1   g731(.A1(new_n869), .A2(new_n610), .A3(new_n927), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n930), .B2(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(G211gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n923), .A2(new_n935), .A3(new_n626), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n869), .A2(new_n626), .A3(new_n926), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n923), .B2(new_n682), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n869), .A2(KEYINPUT126), .A3(new_n927), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(G218gat), .A3(new_n682), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT126), .B1(new_n869), .B2(new_n927), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n943), .B(KEYINPUT127), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1355gat));
endmodule


