//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT65), .B(new_n196), .C1(new_n189), .C2(G137), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n187), .B2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n187), .A2(G134), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n189), .A2(KEYINPUT66), .A3(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n206), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n208), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n213));
  AND4_X1   g027(.A1(new_n198), .A2(new_n204), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n207), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n205), .A2(G143), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n215), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n206), .A3(new_n208), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT11), .B1(new_n187), .B2(G134), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n190), .B(new_n188), .C1(new_n223), .C2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(new_n197), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n226), .B2(new_n198), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT67), .A2(G116), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT67), .A2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n228), .ZN(new_n236));
  OR2_X1    g050(.A1(KEYINPUT67), .A2(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT67), .A2(G116), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(G119), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n214), .A2(new_n227), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G237), .A2(G953), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT27), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n226), .A2(new_n198), .ZN(new_n251));
  INV_X1    g065(.A(new_n222), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n213), .A2(new_n210), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n198), .A3(new_n204), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n216), .A2(new_n215), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n221), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n219), .B2(new_n221), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n204), .A2(new_n210), .A3(new_n213), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(new_n251), .B1(new_n198), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n257), .B(new_n242), .C1(new_n266), .C2(KEYINPUT30), .ZN(new_n267));
  INV_X1    g081(.A(new_n242), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n268), .A3(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n248), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n250), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n250), .A2(new_n267), .A3(KEYINPUT31), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n243), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n268), .B2(new_n266), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n249), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G472), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n284), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n267), .A2(new_n269), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n249), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n291), .B(new_n292), .C1(new_n281), .C2(new_n249), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n268), .B1(new_n253), .B2(new_n256), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n278), .B2(new_n279), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n248), .A2(KEYINPUT29), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n293), .B(new_n285), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G472), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n288), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G221), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n285), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G227), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT75), .ZN(new_n307));
  XNOR2_X1  g121(.A(G110), .B(G140), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n310));
  INV_X1    g124(.A(G104), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(KEYINPUT76), .ZN(new_n312));
  INV_X1    g126(.A(G107), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n312), .A2(new_n314), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(new_n311), .B2(G107), .ZN(new_n320));
  AOI21_X1  g134(.A(G101), .B1(new_n311), .B2(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(G104), .B1(new_n314), .B2(new_n316), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n311), .A2(G107), .ZN(new_n324));
  OAI21_X1  g138(.A(G101), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n322), .A2(new_n325), .A3(new_n210), .A4(new_n213), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n322), .A2(new_n325), .B1(new_n210), .B2(new_n213), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n251), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT12), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n322), .A2(new_n325), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n254), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n326), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n311), .A2(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n319), .A2(new_n320), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n222), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n338), .A2(G101), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(KEYINPUT4), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n251), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n332), .B2(new_n254), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n322), .A4(new_n325), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n309), .B1(new_n336), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n345), .B1(new_n351), .B2(new_n344), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n309), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n309), .ZN(new_n357));
  AOI221_X4 g171(.A(new_n330), .B1(new_n198), .B2(new_n226), .C1(new_n333), .C2(new_n326), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT12), .B1(new_n334), .B2(new_n251), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n349), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n251), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n349), .A3(new_n309), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT78), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n285), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G469), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(G469), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n360), .A2(new_n353), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n309), .B1(new_n364), .B2(new_n349), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n285), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n304), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G217), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(G234), .B2(new_n285), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT22), .B(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n305), .A2(G221), .A3(G234), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n231), .B2(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n231), .A2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G110), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT24), .B(G110), .Z(new_n388));
  XNOR2_X1  g202(.A(G119), .B(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT69), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  INV_X1    g208(.A(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G140), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n396), .A3(KEYINPUT16), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT69), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT16), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n392), .A4(G125), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n205), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n394), .A2(new_n397), .A3(G146), .A4(new_n400), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n391), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G110), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n383), .A2(new_n384), .A3(new_n405), .A4(new_n385), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n389), .B2(new_n388), .ZN(new_n407));
  XNOR2_X1  g221(.A(G125), .B(G140), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n205), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n407), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n381), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n387), .A2(new_n390), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n395), .A2(KEYINPUT16), .A3(G140), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n408), .A2(KEYINPUT16), .B1(new_n413), .B2(new_n398), .ZN(new_n414));
  AOI21_X1  g228(.A(G146), .B1(new_n414), .B2(new_n394), .ZN(new_n415));
  INV_X1    g229(.A(new_n403), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n403), .A3(new_n409), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(KEYINPUT72), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n380), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT72), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n378), .B(new_n379), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT25), .B1(new_n424), .B2(new_n285), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n426));
  NOR4_X1   g240(.A1(new_n420), .A2(new_n423), .A3(new_n426), .A4(G902), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n375), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n404), .A2(new_n410), .A3(new_n381), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n422), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n411), .A2(new_n380), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n285), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n426), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n432), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT73), .A3(new_n375), .ZN(new_n438));
  INV_X1    g252(.A(new_n375), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n285), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT74), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n430), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n305), .A3(G214), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n207), .ZN(new_n448));
  AOI21_X1  g262(.A(G143), .B1(new_n244), .B2(G214), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n207), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n244), .A2(G143), .A3(G214), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n195), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT17), .B(G131), .C1(new_n448), .C2(new_n449), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n402), .A3(new_n403), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT18), .B(G131), .C1(new_n448), .C2(new_n449), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n393), .A2(new_n396), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n462), .A2(new_n409), .A3(KEYINPUT85), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT85), .B1(new_n462), .B2(new_n409), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n459), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G113), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(new_n311), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n457), .A2(new_n465), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  INV_X1    g285(.A(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n450), .A2(new_n454), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n408), .A2(new_n474), .A3(KEYINPUT19), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT19), .B1(new_n408), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n473), .B(new_n403), .C1(new_n477), .C2(G146), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n465), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n469), .A2(new_n471), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT88), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(new_n471), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n472), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  INV_X1    g301(.A(new_n482), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n457), .A2(new_n465), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n472), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n493), .A3(new_n472), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n484), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n285), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n483), .A2(new_n489), .B1(new_n496), .B2(G475), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n209), .A2(G143), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n209), .B2(G143), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n207), .A2(KEYINPUT90), .A3(G128), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(KEYINPUT13), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT13), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n498), .B(new_n502), .C1(new_n503), .C2(KEYINPUT91), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n505), .B(KEYINPUT13), .C1(new_n500), .C2(new_n501), .ZN(new_n506));
  OAI21_X1  g320(.A(G134), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT92), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(G134), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n501), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n189), .A3(new_n498), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n314), .A2(new_n316), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n237), .A2(G122), .A3(new_n238), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n233), .A2(G122), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n510), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT14), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  OAI21_X1  g338(.A(G107), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n511), .A2(new_n189), .A3(new_n498), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n189), .B1(new_n511), .B2(new_n498), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n516), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n302), .A2(new_n374), .A3(G953), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n521), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n521), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n285), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G478), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n535), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G952), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G953), .ZN(new_n541));
  INV_X1    g355(.A(G234), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n446), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n285), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n497), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G214), .B1(G237), .B2(G902), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n338), .A2(G101), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n338), .A2(new_n340), .B1(new_n235), .B2(new_n241), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n332), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n239), .A2(KEYINPUT5), .A3(new_n240), .ZN(new_n556));
  INV_X1    g370(.A(G113), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT5), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n234), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n229), .A2(new_n230), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n234), .B1(new_n560), .B2(G119), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n556), .A2(new_n559), .B1(new_n561), .B2(new_n236), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n565));
  XOR2_X1   g379(.A(G110), .B(G122), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT6), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n552), .A2(new_n553), .B1(new_n555), .B2(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(new_n568), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT80), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n570), .B2(new_n567), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n564), .A2(new_n566), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n213), .A2(new_n395), .A3(new_n210), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n395), .B2(new_n222), .ZN(new_n579));
  INV_X1    g393(.A(G224), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT81), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n579), .B(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n573), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT7), .B1(new_n580), .B2(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n579), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n566), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT83), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n322), .A2(new_n325), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n562), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n562), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n586), .B(new_n592), .C1(new_n564), .C2(new_n566), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(new_n285), .ZN(new_n594));
  OAI21_X1  g408(.A(G210), .B1(G237), .B2(G902), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n584), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n595), .B(KEYINPUT84), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n584), .B2(new_n594), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n550), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n549), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n300), .A2(new_n373), .A3(new_n445), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NOR2_X1   g418(.A1(new_n284), .A2(KEYINPUT93), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n283), .A2(new_n285), .A3(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n274), .A2(new_n275), .B1(new_n281), .B2(new_n249), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n605), .B1(new_n608), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n444), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n595), .B1(new_n584), .B2(new_n594), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n596), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n584), .A2(new_n594), .A3(KEYINPUT94), .A4(new_n595), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n550), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n618), .A3(new_n548), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n533), .B2(new_n534), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(KEYINPUT96), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n521), .A2(new_n531), .ZN(new_n626));
  INV_X1    g440(.A(new_n532), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n521), .A2(new_n531), .A3(new_n532), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n630), .B2(new_n621), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n625), .B1(new_n533), .B2(new_n534), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT33), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n624), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n536), .A2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(G902), .B1(new_n628), .B2(new_n629), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(G478), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n497), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n611), .A2(new_n373), .A3(new_n620), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n538), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n535), .A2(new_n537), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n497), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n611), .A2(new_n373), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n619), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  AND2_X1   g466(.A1(new_n607), .A2(new_n609), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n373), .A2(new_n602), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n417), .A2(new_n418), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n422), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n442), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n430), .A2(new_n438), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n430), .A2(KEYINPUT98), .A3(new_n438), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND4_X1  g481(.A1(new_n300), .A2(new_n373), .A3(new_n662), .A4(new_n663), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n544), .B1(new_n545), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n497), .A2(new_n646), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n596), .A2(new_n614), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n617), .B1(new_n674), .B2(new_n613), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n596), .A2(new_n614), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n550), .B(new_n616), .C1(new_n678), .C2(new_n612), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT99), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n209), .ZN(G30));
  XOR2_X1   g497(.A(new_n670), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n373), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT40), .Z(new_n686));
  OAI21_X1  g500(.A(new_n249), .B1(new_n243), .B2(new_n294), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n272), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n288), .A2(new_n289), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT100), .A4(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n597), .A2(new_n600), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  INV_X1    g510(.A(new_n550), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n489), .A2(new_n483), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n496), .A2(G475), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n646), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n696), .A2(new_n697), .A3(new_n660), .A4(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n686), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NOR2_X1   g518(.A1(new_n668), .A2(new_n679), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n636), .A2(new_n639), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n700), .A4(new_n671), .ZN(new_n708));
  INV_X1    g522(.A(new_n635), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT95), .B1(new_n628), .B2(new_n629), .ZN(new_n710));
  OAI211_X1 g524(.A(KEYINPUT33), .B(new_n632), .C1(new_n710), .C2(new_n625), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(new_n624), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n700), .B(new_n671), .C1(new_n712), .C2(new_n638), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OAI21_X1  g531(.A(new_n700), .B1(new_n712), .B2(new_n638), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n619), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n304), .ZN(new_n720));
  INV_X1    g534(.A(G469), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n357), .B1(new_n352), .B2(new_n361), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n349), .B(new_n309), .C1(new_n358), .C2(new_n359), .ZN(new_n723));
  AOI21_X1  g537(.A(G902), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n372), .B(new_n720), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n370), .A2(new_n371), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n727), .B2(G902), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n720), .A4(new_n372), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n719), .A2(new_n445), .A3(new_n300), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT41), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G113), .ZN(G15));
  NOR2_X1   g548(.A1(new_n619), .A2(new_n647), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n300), .A3(new_n445), .A4(new_n731), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  AND2_X1   g551(.A1(new_n662), .A2(new_n663), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n730), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n739), .A2(new_n549), .A3(new_n679), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n740), .A3(new_n300), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  AOI21_X1  g556(.A(KEYINPUT73), .B1(new_n437), .B2(new_n375), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n429), .B(new_n439), .C1(new_n435), .C2(new_n436), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(G472), .B1(new_n608), .B2(G902), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n284), .A2(new_n285), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n295), .A2(new_n248), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n747), .B1(new_n276), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n443), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n726), .A2(new_n730), .A3(new_n548), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n679), .B2(new_n701), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n698), .A2(new_n699), .B1(new_n645), .B2(new_n644), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n615), .A2(new_n618), .A3(new_n757), .A4(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n754), .A2(new_n759), .A3(KEYINPUT104), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND2_X1  g579(.A1(new_n708), .A2(new_n714), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n283), .A2(new_n285), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n750), .B1(new_n767), .B2(G472), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n731), .A2(new_n675), .A3(new_n660), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT105), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n675), .A2(new_n730), .A3(new_n726), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n660), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n708), .A4(new_n714), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  NAND2_X1  g591(.A1(new_n362), .A2(new_n365), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n721), .B1(new_n778), .B2(new_n285), .ZN(new_n779));
  INV_X1    g593(.A(new_n372), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n720), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n584), .A2(new_n594), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n550), .B(new_n596), .C1(new_n782), .C2(new_n599), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n300), .A2(new_n445), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n715), .A2(new_n785), .A3(KEYINPUT42), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n300), .A2(new_n445), .A3(new_n784), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n766), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND4_X1  g605(.A1(new_n300), .A2(new_n445), .A3(new_n673), .A4(new_n784), .ZN(new_n792));
  XNOR2_X1  g606(.A(KEYINPUT106), .B(G134), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G36));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n355), .B1(new_n350), .B2(new_n354), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n362), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(G469), .B1(new_n778), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT107), .A3(new_n372), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT107), .B1(new_n803), .B2(new_n372), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n720), .B(new_n684), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n712), .A2(new_n638), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n700), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n706), .A2(KEYINPUT43), .A3(new_n497), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(new_n610), .A3(new_n660), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n783), .B1(new_n815), .B2(KEYINPUT44), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n809), .B(new_n816), .C1(KEYINPUT44), .C2(new_n815), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT108), .B(G137), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G39));
  OAI21_X1  g633(.A(new_n720), .B1(new_n806), .B2(new_n807), .ZN(new_n820));
  AND2_X1   g634(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n300), .A2(new_n445), .A3(new_n783), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n715), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n820), .B1(new_n827), .B2(new_n821), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND2_X1  g644(.A1(new_n731), .A2(new_n697), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT116), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n752), .A2(new_n543), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n696), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n783), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n731), .A2(new_n544), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n812), .B2(new_n813), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n660), .A3(new_n768), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n694), .A2(new_n444), .A3(new_n841), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n497), .A3(new_n811), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n728), .A2(new_n372), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n822), .A2(new_n828), .B1(new_n304), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n840), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n846), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n300), .A2(new_n445), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n844), .A2(new_n640), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n834), .A2(new_n675), .A3(new_n731), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n541), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n859), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n852), .B1(new_n846), .B2(new_n851), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n853), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n682), .B1(new_n770), .B2(new_n775), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  INV_X1    g683(.A(new_n781), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n745), .A3(new_n659), .A4(new_n671), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n756), .B2(new_n758), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n705), .A2(new_n715), .B1(new_n694), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n868), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n868), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n754), .A2(new_n759), .A3(KEYINPUT104), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT104), .B1(new_n754), .B2(new_n759), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n741), .A2(new_n732), .A3(new_n736), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT115), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n741), .A2(new_n732), .A3(new_n736), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n764), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n786), .B2(new_n789), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n550), .B(new_n548), .C1(new_n597), .C2(new_n600), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n611), .A2(new_n373), .A3(new_n648), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n664), .B2(new_n654), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(KEYINPUT111), .C1(new_n664), .C2(new_n654), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n611), .A2(new_n373), .A3(new_n640), .A4(new_n891), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n603), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n784), .A2(new_n660), .A3(new_n768), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n792), .B1(new_n766), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n497), .A2(new_n539), .A3(new_n671), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT112), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n903), .A2(new_n783), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n903), .B2(new_n783), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n668), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n889), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n898), .B1(new_n893), .B2(new_n894), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n902), .A2(new_n908), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT114), .A4(new_n896), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n877), .A2(new_n888), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n682), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n872), .A2(new_n694), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n776), .A2(new_n915), .A3(new_n716), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT52), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n868), .A2(new_n873), .A3(new_n869), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n911), .A2(new_n912), .A3(new_n896), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n790), .A2(new_n883), .A3(new_n764), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n886), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n914), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(KEYINPUT53), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n911), .A2(new_n912), .A3(new_n896), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n790), .A2(new_n883), .A3(new_n764), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT53), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n877), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(KEYINPUT54), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n867), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n696), .A2(new_n445), .A3(new_n706), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n847), .A2(KEYINPUT49), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n700), .A2(new_n304), .A3(new_n697), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n694), .B2(new_n939), .ZN(G75));
  NAND2_X1  g754(.A1(new_n540), .A2(G953), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT119), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n914), .A2(new_n923), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(G902), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n599), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n573), .A2(new_n577), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n583), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n942), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n943), .A2(G210), .A3(G902), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(G51));
  INV_X1    g768(.A(new_n942), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT42), .B1(new_n715), .B2(new_n785), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n766), .A2(new_n788), .A3(new_n787), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT53), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n883), .A2(new_n764), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(KEYINPUT115), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n910), .A3(new_n885), .A4(new_n913), .ZN(new_n961));
  INV_X1    g775(.A(new_n876), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n919), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n869), .B1(new_n868), .B2(new_n873), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n965), .A2(new_n927), .A3(new_n928), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT53), .B1(new_n966), .B2(new_n919), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT54), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n925), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n795), .B(KEYINPUT57), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n727), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n944), .A2(new_n798), .A3(new_n800), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n955), .B1(new_n973), .B2(new_n974), .ZN(G54));
  NAND2_X1  g789(.A1(KEYINPUT58), .A2(G475), .ZN(new_n976));
  OR3_X1    g790(.A1(new_n944), .A2(new_n486), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n486), .B1(new_n944), .B2(new_n976), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n955), .B1(new_n977), .B2(new_n978), .ZN(G60));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n932), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT120), .ZN(new_n984));
  INV_X1    g798(.A(new_n634), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n925), .B2(new_n931), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT120), .B1(new_n987), .B2(new_n634), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n985), .A2(new_n981), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n955), .B1(new_n969), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(G63));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  XNOR2_X1  g806(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n374), .A2(new_n285), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n914), .B2(new_n923), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n658), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n942), .B1(new_n997), .B2(new_n424), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n997), .A2(new_n424), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(KEYINPUT61), .A3(new_n942), .A4(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G66));
  INV_X1    g818(.A(new_n546), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n305), .B1(new_n1005), .B2(G224), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n959), .A2(new_n900), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n305), .ZN(new_n1008));
  INV_X1    g822(.A(G898), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n946), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  XOR2_X1   g824(.A(KEYINPUT122), .B(KEYINPUT123), .Z(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1008), .B(new_n1012), .ZN(G69));
  OAI21_X1  g827(.A(new_n257), .B1(new_n266), .B2(KEYINPUT30), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n477), .B(KEYINPUT124), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n868), .A2(new_n716), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n703), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT62), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n685), .A2(new_n783), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1022), .B(new_n854), .C1(new_n640), .C2(new_n648), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n829), .A2(new_n817), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1016), .B1(new_n1026), .B2(new_n305), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1016), .B1(new_n669), .B2(new_n305), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n809), .A2(new_n854), .A3(new_n759), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n817), .A2(new_n790), .A3(new_n792), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n829), .A2(new_n1017), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1028), .B1(new_n1032), .B2(new_n305), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n305), .B1(G227), .B2(G900), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT126), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  OR3_X1    g850(.A1(new_n1027), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1036), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(G72));
  NOR2_X1   g853(.A1(new_n290), .A2(new_n248), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT127), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1030), .A2(new_n1031), .A3(new_n1007), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1045), .B1(new_n291), .B2(new_n272), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n926), .A2(new_n930), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1046), .A2(new_n942), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1044), .B1(new_n1026), .B2(new_n1007), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n249), .B1(new_n267), .B2(new_n269), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G57));
endmodule


