//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n221), .B1(new_n202), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(G77), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G244), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n217), .B2(new_n220), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G222), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G223), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n258), .C1(new_n224), .C2(new_n251), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n209), .A2(new_n262), .B1(new_n216), .B2(new_n256), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n216), .B2(new_n256), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(G226), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT8), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G58), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT68), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n278), .A2(KEYINPUT68), .A3(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n210), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n202), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n275), .B1(G1), .B2(new_n210), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n202), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n272), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n287), .A2(new_n292), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT9), .B1(new_n287), .B2(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n259), .B2(new_n268), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n259), .A2(new_n268), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G190), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n299), .B1(new_n298), .B2(new_n303), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n293), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n251), .A2(new_n315), .A3(G232), .A4(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n251), .A2(G226), .A3(new_n253), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n314), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n258), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n263), .B2(KEYINPUT71), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT71), .B1(new_n257), .B2(new_n266), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n324), .B1(new_n267), .B2(new_n265), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n265), .A2(new_n267), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n257), .A2(new_n266), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT71), .ZN(new_n330));
  OAI21_X1  g0130(.A(G238), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n331), .B2(new_n323), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n258), .B2(new_n319), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n327), .B(G190), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n282), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n273), .A2(new_n274), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n339), .A2(KEYINPUT11), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT12), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n289), .B2(new_n336), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n288), .A2(KEYINPUT12), .A3(G68), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n291), .A2(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n339), .B2(new_n340), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n341), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n335), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n320), .A2(new_n325), .ZN(new_n349));
  INV_X1    g0149(.A(new_n326), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n300), .B1(new_n351), .B2(new_n327), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n308), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n326), .B1(new_n320), .B2(new_n325), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n356), .A2(KEYINPUT73), .A3(new_n347), .A4(new_n335), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n347), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(G169), .C1(new_n354), .C2(new_n355), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n327), .B(G179), .C1(new_n333), .C2(new_n334), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n351), .A2(new_n327), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n360), .B1(new_n364), .B2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n359), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n251), .A2(G232), .A3(new_n253), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n206), .C2(new_n251), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n258), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n263), .A2(new_n225), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n328), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n283), .B1(new_n224), .B2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n277), .A2(new_n279), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n285), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n275), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n291), .A2(new_n338), .B1(new_n224), .B2(new_n288), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(G200), .ZN(new_n385));
  OR3_X1    g0185(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT69), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n374), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G179), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n373), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n372), .B2(new_n271), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n307), .A2(new_n358), .A3(new_n366), .A4(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT77), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n276), .A2(new_n336), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n201), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n285), .A2(KEYINPUT74), .A3(G159), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT74), .B1(new_n285), .B2(G159), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n251), .B2(G20), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n310), .A2(new_n312), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n275), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n311), .B2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n309), .A2(KEYINPUT75), .A3(G33), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n312), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n401), .A2(G20), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n336), .B1(new_n414), .B2(new_n402), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n415), .B2(new_n400), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n280), .A2(new_n281), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n288), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n291), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n407), .A2(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n328), .B1(new_n236), .B2(new_n329), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n251), .A2(new_n427), .A3(G223), .A4(new_n253), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n310), .A2(new_n312), .A3(G223), .A4(new_n253), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n423), .B1(new_n431), .B2(new_n257), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n300), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n423), .B(new_n434), .C1(new_n431), .C2(new_n257), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n421), .A2(new_n436), .A3(KEYINPUT17), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT17), .B1(new_n421), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n394), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n433), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n405), .A2(G68), .ZN(new_n442));
  INV_X1    g0242(.A(new_n400), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT16), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n416), .A3(new_n340), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n420), .A2(new_n418), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n440), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n421), .A2(new_n436), .A3(KEYINPUT17), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT77), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n430), .A2(new_n428), .ZN(new_n451));
  INV_X1    g0251(.A(new_n426), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n257), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G169), .B1(new_n453), .B2(new_n422), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n388), .B2(new_n432), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n447), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n447), .B2(new_n455), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n439), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n273), .A2(new_n274), .B1(G20), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n462), .B2(new_n464), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n288), .A2(G116), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n209), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n275), .A2(new_n288), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(new_n461), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n261), .A2(G1), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n475), .A2(new_n476), .B1(new_n216), .B2(new_n256), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n209), .A2(G45), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n477), .A2(G270), .B1(new_n265), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n309), .A2(G33), .ZN(new_n484));
  OAI21_X1  g0284(.A(G303), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(new_n253), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n310), .A2(new_n312), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n258), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n482), .A2(new_n489), .A3(KEYINPUT82), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n474), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n468), .A2(new_n473), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n482), .A2(new_n489), .A3(G179), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n494), .A2(KEYINPUT21), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n465), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n288), .A2(new_n471), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n340), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n469), .B1(new_n501), .B2(G116), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n271), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n482), .A2(new_n489), .A3(KEYINPUT82), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT82), .B1(new_n482), .B2(new_n489), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n503), .B(KEYINPUT21), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n492), .A2(new_n493), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n503), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n497), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n500), .A2(new_n512), .A3(new_n340), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n376), .A2(new_n288), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n251), .A2(new_n210), .A3(G68), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n210), .B1(new_n317), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G87), .B2(new_n207), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n282), .B2(new_n205), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n513), .B(new_n514), .C1(new_n520), .C2(new_n340), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n257), .A2(G274), .A3(new_n476), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n257), .A2(G250), .A3(new_n478), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n310), .A2(new_n312), .A3(G238), .A4(new_n253), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n528), .B2(new_n258), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n521), .B(new_n530), .C1(new_n300), .C2(new_n529), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n258), .ZN(new_n532));
  INV_X1    g0332(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n271), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n520), .A2(new_n340), .ZN(new_n536));
  INV_X1    g0336(.A(new_n514), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n501), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(new_n388), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n531), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n310), .A2(new_n312), .A3(G250), .A4(new_n253), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G294), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(G1698), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(KEYINPUT87), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n258), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n477), .A2(G264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n481), .A2(new_n265), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n271), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n551), .A3(new_n388), .A4(new_n552), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n310), .A2(new_n312), .A3(new_n210), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n251), .A2(new_n210), .A3(G87), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n206), .A3(G20), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n563), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n556), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n570), .A3(new_n556), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n275), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n288), .B2(G107), .ZN(new_n577));
  AOI22_X1  g0377(.A1(G107), .A2(new_n501), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n554), .B(new_n555), .C1(new_n574), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n553), .A2(G200), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n562), .A2(new_n570), .A3(new_n556), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n340), .B1(new_n582), .B2(new_n571), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n550), .A2(new_n551), .A3(G190), .A4(new_n552), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(new_n583), .A3(new_n578), .A4(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n544), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n504), .B2(new_n505), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n492), .A2(G190), .A3(new_n493), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n495), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT84), .A4(new_n495), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n511), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n477), .A2(G257), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n552), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(new_n253), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(KEYINPUT4), .A2(G244), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n310), .A2(new_n312), .A3(new_n601), .A4(new_n253), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n463), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n310), .A2(new_n312), .A3(G250), .A4(G1698), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n251), .A2(KEYINPUT78), .A3(G250), .A4(G1698), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n258), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n258), .C1(new_n603), .C2(new_n608), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n597), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n595), .B1(new_n613), .B2(new_n300), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n596), .A2(new_n552), .ZN(new_n615));
  INV_X1    g0415(.A(new_n612), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n602), .A2(new_n463), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n600), .A3(new_n606), .A4(new_n607), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n611), .B1(new_n618), .B2(new_n258), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(KEYINPUT80), .A3(G200), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n285), .A2(G77), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT6), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n623), .A2(new_n205), .A3(G107), .ZN(new_n624));
  XNOR2_X1  g0424(.A(G97), .B(G107), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(new_n210), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n206), .B1(new_n414), .B2(new_n402), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n340), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n288), .A2(G97), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n501), .B2(G97), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n609), .A2(new_n615), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n629), .B(new_n631), .C1(new_n632), .C2(new_n434), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n614), .A2(new_n621), .A3(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n388), .B(new_n615), .C1(new_n616), .C2(new_n619), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n632), .A2(new_n271), .B1(new_n629), .B2(new_n631), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NOR4_X1   g0439(.A1(new_n393), .A2(new_n460), .A3(new_n594), .A4(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n293), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n356), .A2(new_n347), .A3(new_n335), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n389), .A3(new_n390), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n366), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT90), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n366), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n645), .A2(new_n439), .A3(new_n450), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n459), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n304), .A2(new_n305), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n641), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n393), .A2(new_n460), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n508), .A2(new_n510), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n495), .A2(new_n496), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n509), .A2(new_n503), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(new_n657), .A3(new_n580), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n534), .A2(KEYINPUT88), .A3(G200), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n529), .B2(new_n300), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(new_n661), .A3(new_n530), .A4(new_n521), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n585), .A2(new_n543), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n658), .A2(new_n638), .A3(new_n635), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(new_n638), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n544), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n543), .B(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n636), .A2(new_n637), .A3(new_n662), .A4(new_n543), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n652), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n651), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n653), .A2(new_n657), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n591), .B2(new_n592), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n495), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g0485(.A(new_n677), .B(new_n676), .S(new_n685), .Z(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n580), .A2(new_n683), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n683), .B1(new_n574), .B2(new_n579), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n585), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n691), .B2(new_n580), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n689), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n676), .A2(new_n684), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n692), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n694), .A3(new_n698), .ZN(G399));
  NAND2_X1  g0499(.A1(new_n213), .A2(new_n260), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT92), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n220), .B2(new_n700), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n703), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n609), .A2(new_n615), .A3(new_n551), .A4(new_n550), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n529), .A2(G179), .A3(new_n482), .A4(new_n489), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT30), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n496), .A2(new_n534), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n550), .A2(new_n551), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n597), .B1(new_n618), .B2(new_n258), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n529), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n620), .A2(new_n509), .A3(new_n553), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n683), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n684), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n723), .A2(new_n724), .B1(new_n719), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n639), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n677), .A2(new_n727), .A3(new_n586), .A4(new_n684), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n707), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n635), .A2(new_n663), .A3(new_n638), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n653), .A2(new_n657), .A3(new_n580), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n666), .A2(new_n665), .A3(new_n544), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n670), .A2(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n669), .A3(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT29), .B(new_n684), .C1(new_n733), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n683), .B1(new_n664), .B2(new_n672), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(KEYINPUT29), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n706), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(new_n700), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n210), .A2(G13), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n209), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n743), .A2(KEYINPUT94), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT94), .B1(new_n743), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n688), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n686), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n274), .B1(G20), .B2(new_n271), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(G190), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n388), .A3(new_n300), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G159), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n757), .A2(new_n758), .B1(new_n336), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n757), .B2(new_n758), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n210), .A2(new_n434), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n388), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n251), .B1(new_n766), .B2(new_n276), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n754), .A2(new_n765), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(new_n224), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n434), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n210), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n205), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n759), .A2(new_n434), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(G50), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT97), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n300), .B2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n388), .A2(KEYINPUT97), .A3(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n778), .A3(new_n754), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G87), .A2(new_n780), .B1(new_n782), .B2(G107), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n763), .A2(new_n770), .A3(new_n775), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n772), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(KEYINPUT33), .A2(G317), .ZN(new_n787));
  NAND2_X1  g0587(.A1(KEYINPUT33), .A2(G317), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n761), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n786), .B(new_n789), .C1(G326), .C2(new_n774), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n782), .A2(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n768), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n403), .B1(new_n766), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G329), .C2(new_n756), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n780), .A2(G303), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n790), .A2(new_n791), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n784), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n753), .B1(new_n800), .B2(KEYINPUT98), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(KEYINPUT98), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n213), .A2(new_n251), .ZN(new_n803));
  INV_X1    g0603(.A(G355), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(G116), .B2(new_n213), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n246), .A2(new_n261), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT95), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n213), .A2(new_n403), .ZN(new_n808));
  INV_X1    g0608(.A(new_n220), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n261), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n805), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n753), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n750), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n802), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n814), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n686), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n752), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NOR2_X1   g0622(.A1(new_n391), .A2(new_n683), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n387), .B1(new_n382), .B2(new_n684), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n391), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n738), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n749), .B1(new_n826), .B2(new_n730), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(KEYINPUT101), .B1(new_n730), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(KEYINPUT101), .B2(new_n828), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n403), .B1(new_n756), .B2(G132), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n782), .A2(G68), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n276), .C2(new_n772), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G137), .A2(new_n774), .B1(new_n760), .B2(G150), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT100), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  INV_X1    g0636(.A(G159), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n766), .C1(new_n837), .C2(new_n768), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  AOI211_X1 g0639(.A(new_n833), .B(new_n839), .C1(G50), .C2(new_n780), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n403), .B1(new_n766), .B2(new_n785), .C1(new_n792), .C2(new_n755), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n773), .B(new_n841), .C1(G303), .C2(new_n774), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n842), .B1(new_n512), .B2(new_n781), .C1(new_n206), .C2(new_n779), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n761), .A2(new_n844), .B1(new_n768), .B2(new_n461), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n753), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n753), .A2(new_n812), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n749), .B1(new_n338), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(new_n813), .C2(new_n825), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n830), .A2(new_n851), .ZN(G384));
  OAI211_X1 g0652(.A(new_n737), .B(new_n652), .C1(KEYINPUT29), .C2(new_n738), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n651), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT106), .Z(new_n855));
  NAND2_X1  g0655(.A1(new_n444), .A2(new_n340), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n446), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n681), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n460), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n455), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n421), .A2(new_n436), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n447), .A2(new_n455), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n447), .A2(new_n859), .ZN(new_n868));
  XOR2_X1   g0668(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n869));
  NAND4_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  AOI221_X4 g0677(.A(new_n873), .B1(new_n866), .B2(new_n870), .C1(new_n460), .C2(new_n861), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n437), .A2(new_n438), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n868), .B1(new_n459), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n867), .A2(new_n868), .A3(new_n864), .ZN(new_n882));
  INV_X1    g0682(.A(new_n869), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n870), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n877), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n876), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(G169), .B1(new_n354), .B2(new_n355), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT14), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n362), .A3(new_n361), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n359), .A3(new_n684), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n874), .A2(new_n875), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n738), .A2(new_n825), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n823), .B(KEYINPUT103), .Z(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n347), .A2(new_n684), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n642), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n366), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n363), .A2(new_n365), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n358), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  AOI211_X1 g0708(.A(KEYINPUT104), .B(new_n902), .C1(new_n358), .C2(new_n906), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n896), .A2(new_n900), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n459), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n681), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n895), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n855), .B(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n825), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n892), .B1(new_n353), .B2(new_n357), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT104), .B1(new_n917), .B2(new_n902), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n907), .A2(new_n905), .A3(new_n901), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n920), .B2(new_n904), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n553), .B(new_n717), .C1(new_n504), .C2(new_n505), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n620), .A2(new_n923), .B1(new_n710), .B2(new_n715), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n683), .B1(new_n924), .B2(new_n721), .ZN(new_n925));
  INV_X1    g0725(.A(new_n722), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n724), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n683), .A4(new_n722), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n728), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n921), .B(new_n929), .C1(new_n878), .C2(new_n886), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT40), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n896), .A2(new_n921), .A3(new_n932), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n652), .ZN(new_n936));
  OAI21_X1  g0736(.A(G330), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n915), .A2(new_n938), .B1(new_n209), .B2(new_n744), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n915), .B2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n626), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n942), .A2(G20), .A3(G116), .A4(new_n216), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT102), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n943), .A2(new_n944), .B1(new_n941), .B2(new_n626), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n809), .B(new_n224), .C1(new_n276), .C2(new_n336), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n202), .A2(G68), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n209), .B(G13), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n940), .A2(new_n947), .A3(new_n950), .ZN(G367));
  AOI21_X1  g0751(.A(new_n684), .B1(new_n629), .B2(new_n631), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n639), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n666), .A2(new_n683), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n698), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n638), .B1(new_n953), .B2(new_n580), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n684), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n662), .A2(new_n543), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n521), .A2(new_n684), .ZN(new_n962));
  MUX2_X1   g0762(.A(new_n961), .B(new_n669), .S(new_n962), .Z(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n960), .A2(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n693), .A2(new_n955), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n967), .C1(new_n970), .C2(new_n971), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n700), .B(KEYINPUT41), .ZN(new_n977));
  INV_X1    g0777(.A(new_n955), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n698), .A3(new_n694), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n698), .B2(new_n694), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n693), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n697), .B(new_n692), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n688), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n741), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n980), .A2(new_n982), .A3(new_n693), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n977), .B1(new_n990), .B2(new_n741), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT108), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n745), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g0793(.A(KEYINPUT108), .B(new_n977), .C1(new_n990), .C2(new_n741), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n975), .B(new_n976), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G150), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n766), .A2(new_n996), .B1(new_n768), .B2(new_n202), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n403), .B(new_n997), .C1(G137), .C2(new_n756), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n780), .A2(G58), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n782), .A2(new_n224), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n772), .A2(new_n336), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n774), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n837), .B2(new_n761), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n779), .A2(new_n461), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT46), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n772), .A2(new_n206), .B1(new_n761), .B2(new_n785), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G311), .B2(new_n774), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n782), .A2(G97), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT109), .B(G317), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n251), .B1(new_n756), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n766), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G303), .A2(new_n1012), .B1(new_n769), .B2(G283), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1001), .A2(new_n1004), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n753), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n815), .B1(new_n213), .B2(new_n375), .C1(new_n242), .C2(new_n808), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n750), .A3(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n963), .A2(new_n814), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n1022), .ZN(G387));
  OR2_X1    g0823(.A1(new_n692), .A2(new_n819), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n803), .A2(new_n701), .B1(G107), .B2(new_n213), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n239), .A2(new_n261), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n701), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1027), .C1(G68), .C2(G77), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n378), .A2(new_n202), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT50), .Z(new_n1030));
  AOI21_X1  g0830(.A(new_n808), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1025), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n750), .B1(new_n1032), .B2(new_n816), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n251), .B1(new_n755), .B2(new_n996), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n766), .A2(new_n202), .B1(new_n768), .B2(new_n336), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G159), .C2(new_n774), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n538), .A2(new_n539), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n772), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n419), .A2(new_n760), .B1(new_n780), .B2(new_n224), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1009), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1012), .A2(new_n1010), .B1(new_n769), .B2(G303), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n774), .A2(G322), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n792), .C2(new_n761), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n844), .A2(new_n772), .B1(new_n779), .B2(new_n785), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n251), .B1(new_n756), .B2(G326), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n461), .C2(new_n781), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1041), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n1053), .B2(new_n753), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n986), .A2(new_n746), .B1(new_n1024), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n700), .B(KEYINPUT110), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n987), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n986), .A2(new_n741), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(G393));
  NAND2_X1  g0859(.A1(new_n990), .A2(new_n1056), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n989), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT111), .B1(new_n1061), .B2(new_n983), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n983), .A2(KEYINPUT111), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(new_n1064), .B2(new_n987), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n815), .B1(new_n205), .B2(new_n213), .C1(new_n249), .C2(new_n808), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n750), .A2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1012), .A2(G311), .B1(G317), .B2(new_n774), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n403), .B1(new_n768), .B2(new_n785), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G322), .B2(new_n756), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1038), .A2(G116), .B1(G303), .B2(new_n760), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G283), .A2(new_n780), .B1(new_n782), .B2(G107), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT112), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1012), .A2(G159), .B1(G150), .B2(new_n774), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  AOI21_X1  g0878(.A(new_n403), .B1(new_n769), .B2(new_n378), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n836), .B2(new_n755), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n772), .A2(new_n338), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G50), .B2(new_n760), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G68), .A2(new_n780), .B1(new_n782), .B2(G87), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1078), .A2(new_n1081), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1076), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1067), .B1(new_n1087), .B2(new_n753), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n978), .B2(new_n819), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1064), .B2(new_n745), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1065), .A2(new_n1090), .ZN(G390));
  AOI21_X1  g0891(.A(new_n898), .B1(new_n738), .B2(new_n825), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n918), .A2(new_n919), .B1(new_n366), .B2(new_n903), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n893), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n684), .B1(new_n733), .B2(new_n736), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n899), .B1(new_n1095), .B2(new_n916), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n910), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n885), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n873), .B1(new_n1098), .B2(new_n880), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n894), .B1(new_n875), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n888), .A2(new_n1094), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n910), .A2(new_n929), .A3(G330), .A4(new_n825), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT113), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n729), .A2(new_n910), .A3(new_n825), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT114), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n921), .A2(new_n1106), .A3(new_n729), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1102), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n900), .A2(new_n910), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n893), .B1(new_n876), .B2(new_n887), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1110), .B(new_n1111), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1103), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n746), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n849), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n750), .B1(new_n419), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n755), .A2(new_n785), .B1(new_n768), .B2(new_n205), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n251), .B(new_n1120), .C1(G116), .C2(new_n1012), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n780), .A2(G87), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n832), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1082), .B1(G283), .B2(new_n774), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n206), .B2(new_n761), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n780), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n760), .A2(G137), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n772), .B2(new_n837), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n774), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n782), .A2(G50), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n403), .B1(new_n769), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G125), .A2(new_n756), .B1(new_n1012), .B2(G132), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1123), .A2(new_n1125), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1119), .B1(new_n1136), .B2(new_n753), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n889), .B2(new_n813), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n719), .A2(new_n725), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n927), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n594), .A2(new_n639), .A3(new_n683), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n825), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1093), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1092), .B1(new_n1144), .B2(new_n1102), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n929), .A2(G330), .A3(new_n825), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1096), .B1(new_n1146), .B2(new_n1093), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1108), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n366), .A2(new_n646), .A3(new_n643), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n646), .B1(new_n366), .B2(new_n643), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n439), .A2(new_n450), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n650), .B1(new_n1152), .B2(new_n912), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n927), .A2(new_n928), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n652), .C1(new_n1154), .C2(new_n1142), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n853), .A2(new_n1153), .A3(new_n1155), .A4(new_n293), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT115), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n651), .A2(KEYINPUT115), .A3(new_n853), .A4(new_n1155), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1139), .B1(new_n1148), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n921), .A2(new_n1106), .A3(new_n729), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1106), .B1(new_n921), .B2(new_n729), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1147), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1145), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT116), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1169), .A2(KEYINPUT117), .A3(new_n1116), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT117), .B1(new_n1169), .B2(new_n1116), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1056), .B1(new_n1169), .B2(new_n1116), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1117), .B(new_n1138), .C1(new_n1172), .C2(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n934), .A2(G330), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1176));
  OR2_X1    g0976(.A1(new_n306), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n294), .A2(new_n681), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n306), .A2(new_n1176), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1179), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1175), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n914), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1183), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n934), .A2(new_n1186), .A3(G330), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n934), .B2(G330), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n707), .B(new_n1183), .C1(new_n931), .C2(new_n933), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n914), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1191), .A3(KEYINPUT121), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n914), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT121), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1183), .A2(new_n812), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n750), .B1(G50), .B2(new_n1118), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n780), .A2(new_n224), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n756), .A2(G283), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1012), .A2(G107), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n251), .A2(G41), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1037), .B2(new_n769), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n782), .A2(G58), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT118), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n761), .A2(new_n205), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1207), .B(new_n1002), .C1(G116), .C2(new_n774), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1202), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1038), .A2(G150), .B1(G125), .B2(new_n774), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G128), .A2(new_n1012), .B1(new_n769), .B2(G137), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n780), .A2(new_n1132), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n760), .A2(G132), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n782), .A2(G159), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n756), .C2(G124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1214), .B1(new_n1210), .B2(new_n1209), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1198), .B1(new_n1225), .B2(new_n753), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1196), .A2(new_n746), .B1(new_n1197), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1169), .A2(new_n1116), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT117), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1169), .A2(KEYINPUT117), .A3(new_n1116), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1160), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1191), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1193), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1056), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1196), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1227), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT122), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1240), .B(new_n1227), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n1093), .A2(new_n812), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n749), .B1(new_n336), .B2(new_n849), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1039), .B1(new_n338), .B2(new_n781), .C1(new_n205), .C2(new_n779), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G283), .A2(new_n1012), .B1(new_n769), .B2(G107), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n251), .B1(new_n756), .B2(G303), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G116), .A2(new_n760), .B1(new_n774), .B2(G294), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1132), .A2(new_n760), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n202), .B2(new_n772), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G132), .B2(new_n774), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n780), .A2(G159), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n403), .B1(new_n769), .B2(G150), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G128), .A2(new_n756), .B1(new_n1012), .B2(G137), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1206), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1247), .A2(new_n1251), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1246), .B1(new_n753), .B2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1166), .A2(new_n746), .B1(new_n1244), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1148), .A2(new_n1160), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT123), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1169), .A2(new_n977), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1263), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(G381));
  OR4_X1    g1069(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1270), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1242), .ZN(G407));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(G378), .A2(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1242), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1273), .B1(new_n1242), .B2(new_n1277), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(new_n1278), .C2(new_n1279), .ZN(G409));
  INV_X1    g1080(.A(G390), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n975), .A2(new_n976), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n990), .A2(new_n741), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n977), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n746), .B1(new_n1285), .B2(KEYINPUT108), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n994), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1282), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1281), .B1(new_n1288), .B2(new_n1021), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n995), .A2(G390), .A3(new_n1022), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(G393), .B(new_n821), .ZN(new_n1291));
  AND4_X1   g1091(.A1(KEYINPUT127), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1294), .A2(new_n1291), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1227), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1117), .A2(new_n1138), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1172), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1173), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1236), .A2(new_n1284), .A3(new_n1196), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n746), .B1(new_n1233), .B2(new_n1193), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1197), .A2(new_n1226), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1276), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1161), .A2(new_n1168), .A3(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1266), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1056), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1313), .B1(new_n1264), .B2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1148), .A2(KEYINPUT126), .A3(KEYINPUT60), .A4(new_n1160), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1312), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1311), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1318), .B2(new_n1262), .ZN(new_n1319));
  INV_X1    g1119(.A(G384), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1320), .B(new_n1263), .C1(new_n1311), .C2(new_n1317), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1297), .B1(new_n1309), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1262), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1320), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1318), .A2(G384), .A3(new_n1262), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1275), .A2(G2897), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1328), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1330), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1275), .B1(new_n1298), .B2(new_n1307), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1322), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1296), .A2(new_n1324), .A3(new_n1333), .A4(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1334), .A2(new_n1337), .A3(new_n1322), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1339), .B1(new_n1334), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1337), .B1(new_n1334), .B2(new_n1322), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1338), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1336), .B1(new_n1343), .B2(new_n1296), .ZN(G405));
  NAND3_X1  g1144(.A1(new_n1239), .A2(new_n1302), .A3(new_n1241), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1323), .A3(new_n1298), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1323), .B1(new_n1345), .B2(new_n1298), .ZN(new_n1348));
  OAI22_X1  g1148(.A1(new_n1347), .A2(new_n1348), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1348), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1296), .A3(new_n1346), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(G402));
endmodule


