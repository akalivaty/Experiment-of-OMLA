//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT67), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G238), .A2(G237), .A3(G236), .A4(G235), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT69), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT70), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n459), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n459), .B1(new_n465), .B2(new_n467), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT71), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n484), .B2(G124), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n462), .A2(new_n468), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n464), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(KEYINPUT72), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n459), .B2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n493), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n489), .A2(new_n486), .A3(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n483), .A2(G126), .B1(new_n473), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n490), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND4_X1   g091(.A1(new_n506), .A2(new_n508), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n514), .A2(new_n516), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n513), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G543), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n517), .A2(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(new_n509), .A2(new_n520), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n509), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n504), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n506), .A2(new_n508), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n504), .B1(new_n546), .B2(KEYINPUT75), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(KEYINPUT75), .B2(new_n546), .ZN(new_n548));
  INV_X1    g123(.A(new_n531), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G43), .B1(G81), .B2(new_n517), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n544), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT78), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G65), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(KEYINPUT79), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G651), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n564), .A2(KEYINPUT80), .A3(G651), .A4(new_n565), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n520), .A2(KEYINPUT77), .A3(G53), .A4(G543), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n572), .B(KEYINPUT9), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n517), .A2(G91), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n568), .A2(new_n569), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n582));
  INV_X1    g157(.A(new_n524), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(new_n522), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n584), .B2(new_n513), .ZN(new_n585));
  AOI211_X1 g160(.A(KEYINPUT81), .B(new_n512), .C1(new_n583), .C2(new_n522), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G303));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  INV_X1    g163(.A(G49), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n535), .A2(new_n588), .B1(new_n531), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n549), .A2(G48), .B1(G86), .B2(new_n517), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n504), .B2(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n504), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n549), .A2(G47), .B1(G85), .B2(new_n517), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n558), .A2(new_n559), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n504), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n535), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n612), .A2(new_n613), .B1(G54), .B2(new_n549), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(new_n551), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n619), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n615), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g204(.A1(new_n462), .A2(new_n468), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n630), .A2(G2104), .A3(new_n459), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n484), .A2(G123), .ZN(new_n637));
  INV_X1    g212(.A(new_n478), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n637), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n636), .A3(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(KEYINPUT17), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(new_n668), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n662), .B(new_n669), .S(new_n673), .Z(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT20), .Z(new_n688));
  OR2_X1    g263(.A1(new_n681), .A2(new_n683), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n686), .A3(new_n684), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n688), .B(new_n690), .C1(new_n686), .C2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT86), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G20), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT94), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT23), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G299), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT95), .ZN(new_n704));
  INV_X1    g279(.A(G1956), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g284(.A(G140), .ZN(new_n710));
  NOR2_X1   g285(.A1(G104), .A2(G2105), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n478), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n484), .B2(G128), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2067), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT25), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n630), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n459), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n718), .B(new_n720), .C1(G139), .C2(new_n638), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n707), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n707), .B2(G33), .ZN(new_n723));
  INV_X1    g298(.A(G2072), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  INV_X1    g300(.A(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G160), .B2(new_n707), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n723), .A2(new_n724), .B1(G2084), .B2(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n716), .B(new_n730), .C1(new_n724), .C2(new_n723), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n699), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n699), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1961), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n707), .A2(G32), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G141), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n478), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G129), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n734), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n707), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n748), .B1(new_n750), .B2(new_n751), .C1(new_n642), .C2(new_n707), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n699), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n699), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n752), .B1(new_n754), .B2(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n707), .A2(G27), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G164), .B2(new_n707), .ZN(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n729), .A2(G2084), .ZN(new_n760));
  AND4_X1   g335(.A1(new_n746), .A2(new_n755), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n699), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n616), .B2(new_n699), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT91), .B(G1348), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G19), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n551), .B2(new_n699), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1341), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n731), .A2(new_n761), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n707), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n707), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT29), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n754), .A2(G1966), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n744), .A2(new_n745), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n776), .B(new_n777), .C1(G1961), .C2(new_n733), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n773), .A2(new_n774), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR4_X1    g355(.A1(new_n706), .A2(new_n770), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  MUX2_X1   g357(.A(G6), .B(G305), .S(G16), .Z(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT89), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT90), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n699), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n699), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1971), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n699), .A2(G23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n593), .B2(new_n699), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n787), .A2(new_n788), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n798));
  INV_X1    g373(.A(G25), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n799), .A2(KEYINPUT87), .A3(G29), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT87), .B1(new_n799), .B2(G29), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G107), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n464), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n638), .A2(G131), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n484), .B2(G119), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n800), .B(new_n801), .C1(new_n807), .C2(new_n707), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n699), .A2(G24), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT88), .Z(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n699), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n810), .B1(new_n814), .B2(G1986), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G1986), .B2(new_n814), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n797), .A2(new_n798), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT36), .Z(new_n818));
  NOR2_X1   g393(.A1(new_n782), .A2(new_n818), .ZN(G311));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n781), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(G150));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n535), .A2(new_n824), .B1(new_n531), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT97), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(new_n504), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n616), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT38), .Z(new_n835));
  AND2_X1   g410(.A1(new_n827), .A2(new_n829), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n625), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n551), .A3(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n835), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n833), .B1(new_n846), .B2(new_n848), .ZN(G145));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  NOR2_X1   g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n478), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n484), .B2(G130), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n632), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n807), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT100), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n714), .B(new_n502), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n743), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n721), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n642), .B(G160), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n856), .ZN(new_n865));
  INV_X1    g440(.A(new_n863), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n865), .B(new_n866), .C1(new_n857), .C2(new_n860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g444(.A(new_n843), .B(new_n627), .ZN(new_n870));
  XNOR2_X1  g445(.A(G299), .B(new_n616), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G299), .B(new_n615), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n871), .B2(new_n870), .ZN(new_n879));
  XNOR2_X1  g454(.A(G290), .B(G166), .ZN(new_n880));
  XNOR2_X1  g455(.A(G288), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT42), .Z(new_n883));
  OR2_X1    g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n619), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n836), .A2(G868), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n886), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT101), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(G295));
  OR2_X1    g465(.A1(new_n886), .A2(new_n887), .ZN(G331));
  XNOR2_X1  g466(.A(G168), .B(G171), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n842), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n551), .B1(new_n838), .B2(new_n839), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n841), .A2(new_n842), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n876), .ZN(new_n899));
  INV_X1    g474(.A(new_n882), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n871), .A3(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n905), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n905), .B2(G37), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n906), .B2(new_n902), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n912), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n904), .ZN(new_n918));
  MUX2_X1   g493(.A(new_n915), .B(new_n918), .S(KEYINPUT44), .Z(G397));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n488), .A2(new_n489), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n473), .A2(new_n500), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT72), .B1(new_n492), .B2(new_n494), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n497), .A2(new_n496), .A3(new_n493), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n920), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G160), .A2(G40), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(G1996), .A3(new_n743), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT103), .Z(new_n933));
  XNOR2_X1  g508(.A(new_n714), .B(G2067), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G1996), .B2(new_n743), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n807), .B(new_n809), .Z(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n525), .A2(KEYINPUT81), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n584), .A2(new_n582), .A3(new_n513), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(G8), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT55), .A4(G8), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n920), .ZN(new_n954));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n472), .A2(new_n955), .A3(new_n476), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT45), .B1(new_n502), .B2(new_n920), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n929), .A2(new_n960), .A3(new_n956), .A4(new_n954), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT105), .B(G1971), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n930), .B1(KEYINPUT50), .B2(new_n927), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n927), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n502), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(G2090), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n953), .A2(G8), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(G8), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n502), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT106), .B1(new_n502), .B2(new_n920), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n977), .B2(new_n956), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n593), .A2(G1976), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT109), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n966), .A2(new_n956), .A3(new_n968), .ZN(new_n983));
  INV_X1    g558(.A(new_n974), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n979), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(KEYINPUT109), .B2(new_n980), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n593), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(G305), .A2(G1981), .ZN(new_n989));
  NOR2_X1   g564(.A1(G305), .A2(G1981), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n978), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n990), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n978), .B(KEYINPUT110), .Z(new_n998));
  OAI22_X1  g573(.A1(new_n973), .A2(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g576(.A(G1966), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n966), .B2(new_n968), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n957), .ZN(new_n1004));
  INV_X1    g579(.A(G2084), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n964), .A2(new_n969), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G168), .A2(new_n974), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT122), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT122), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g592(.A(KEYINPUT51), .B(new_n1008), .C1(new_n1007), .C2(new_n984), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1001), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1016), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1008), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1015), .B2(KEYINPUT122), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT62), .B(new_n1020), .C1(new_n1024), .C2(new_n1010), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1003), .ZN(new_n1026));
  INV_X1    g601(.A(new_n957), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n758), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1961), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n970), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G2078), .B1(new_n959), .B2(new_n961), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1028), .B(new_n1030), .C1(new_n1031), .C2(KEYINPUT53), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G301), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1019), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n953), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n967), .B1(new_n966), .B2(new_n968), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n930), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT111), .B(new_n956), .C1(new_n977), .C2(new_n967), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n502), .A2(new_n967), .A3(new_n920), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n774), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n963), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT112), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n984), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(KEYINPUT112), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n988), .A2(new_n1049), .A3(new_n994), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n972), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1000), .B1(new_n1035), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n705), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n957), .A2(new_n958), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G299), .A2(KEYINPUT115), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n566), .B2(new_n567), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n569), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1060), .A2(new_n1064), .A3(KEYINPUT57), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n970), .A2(new_n764), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n983), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n966), .A2(KEYINPUT116), .A3(new_n956), .A4(new_n968), .ZN(new_n1073));
  AOI21_X1  g648(.A(G2067), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT117), .B(G2067), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2067), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n977), .B2(new_n956), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1073), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(KEYINPUT118), .A3(new_n1084), .A4(new_n1070), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1085), .A3(new_n616), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1068), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1078), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n615), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n616), .A2(KEYINPUT121), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1093), .B(new_n1095), .C1(new_n1078), .C2(new_n1085), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(G1341), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1072), .A2(new_n1073), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1996), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1102), .A2(new_n1103), .B1(new_n1105), .B2(new_n1056), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n551), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1110), .A3(new_n551), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1060), .A2(new_n1064), .A3(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1054), .A2(new_n705), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1087), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1087), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1112), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1089), .B1(new_n1099), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n958), .A2(new_n930), .A3(KEYINPUT123), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n929), .B2(new_n956), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n954), .A2(KEYINPUT53), .A3(new_n758), .ZN(new_n1130));
  OAI221_X1 g705(.A(new_n1030), .B1(new_n1129), .B2(new_n1130), .C1(new_n1031), .C2(KEYINPUT53), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1131), .B2(G171), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1033), .A2(G301), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT124), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1131), .A2(G171), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1125), .B1(new_n1034), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1136), .A2(new_n1047), .A3(new_n1051), .A4(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1053), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1007), .A2(new_n984), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G286), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1047), .A2(new_n1051), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT114), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(KEYINPUT114), .A3(new_n1145), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n973), .A2(KEYINPUT63), .A3(new_n1143), .ZN(new_n1149));
  INV_X1    g724(.A(new_n995), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n971), .A2(G8), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n953), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1147), .A2(new_n1148), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n943), .B1(new_n1141), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n941), .A2(new_n931), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT48), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n939), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT46), .ZN(new_n1160));
  INV_X1    g735(.A(new_n931), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(G1996), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n931), .A2(KEYINPUT46), .A3(new_n1105), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n934), .A2(new_n742), .A3(new_n741), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1162), .B(new_n1163), .C1(new_n1164), .C2(new_n1161), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1166));
  XNOR2_X1  g741(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n809), .B(new_n806), .C1(G119), .C2(new_n484), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n936), .A2(new_n1169), .B1(new_n1079), .B2(new_n714), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1161), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n1156), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n943), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1019), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n999), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1095), .B1(new_n1179), .B2(new_n1093), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1091), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT61), .B1(new_n1068), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1087), .A2(new_n1120), .A3(new_n1113), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1184), .A2(new_n1185), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1088), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1134), .B(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1189), .A2(new_n1177), .A3(new_n1138), .A4(new_n1136), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1178), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1144), .A2(KEYINPUT114), .A3(new_n1145), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1192), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1175), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(new_n1172), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1174), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g772(.A1(new_n677), .A2(G319), .A3(new_n660), .A4(new_n678), .ZN(new_n1199));
  AOI211_X1 g773(.A(new_n1199), .B(G229), .C1(new_n864), .C2(new_n867), .ZN(new_n1200));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n1200), .A2(new_n915), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1201), .B1(new_n1200), .B2(new_n915), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n915), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1205), .A2(KEYINPUT127), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n1200), .A2(new_n915), .A3(new_n1201), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1207), .ZN(G225));
endmodule


