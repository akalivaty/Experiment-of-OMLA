//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1265, new_n1266, new_n1267, new_n1268;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n466), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n462), .A2(G136), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n460), .B2(new_n461), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G162));
  OAI21_X1  g052(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n480), .B2(G114), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT69), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n463), .C1(new_n485), .C2(new_n486), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G138), .A4(new_n463), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n489), .A2(new_n491), .B1(new_n493), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI211_X1 g083(.A(G88), .B(new_n501), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(G50), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(new_n506), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n501), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT72), .Z(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n498), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT71), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n509), .B2(new_n510), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n498), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  INV_X1    g104(.A(new_n501), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n531));
  INV_X1    g106(.A(new_n508), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n529), .B1(new_n533), .B2(G89), .ZN(new_n534));
  OAI211_X1 g109(.A(G51), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT74), .B1(new_n535), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(KEYINPUT75), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n533), .A2(G90), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n531), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G52), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(G651), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n547), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  OAI21_X1  g127(.A(new_n532), .B1(new_n549), .B2(new_n502), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n553), .A2(G81), .A3(new_n501), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(G43), .A3(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n499), .B2(new_n500), .ZN(new_n557));
  AND2_X1   g132(.A1(G68), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n516), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT76), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n554), .A2(new_n555), .A3(new_n562), .A4(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  OAI211_X1 g145(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n553), .A2(new_n573), .A3(G53), .A4(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n508), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n576), .B2(new_n530), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n553), .A2(new_n578), .A3(new_n501), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(G91), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n503), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n575), .A2(new_n580), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  NAND3_X1  g159(.A1(new_n577), .A2(G87), .A3(new_n579), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n503), .B1(new_n530), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n546), .B2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n501), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n549), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(G48), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n553), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n577), .A2(G86), .A3(new_n579), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  XNOR2_X1  g171(.A(KEYINPUT78), .B(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n533), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n546), .A2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n549), .C2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n577), .A2(G92), .A3(new_n579), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n579), .A4(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n546), .A2(G54), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n503), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n612), .B1(new_n606), .B2(new_n607), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n603), .B1(new_n619), .B2(new_n602), .ZN(G321));
  XNOR2_X1  g195(.A(G321), .B(KEYINPUT80), .ZN(G284));
  XNOR2_X1  g196(.A(G299), .B(KEYINPUT81), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n622), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XOR2_X1   g199(.A(KEYINPUT83), .B(G559), .Z(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(G860), .B2(new_n625), .ZN(G148));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n602), .B1(new_n619), .B2(new_n625), .ZN(new_n628));
  AOI211_X1 g203(.A(new_n627), .B(new_n628), .C1(new_n602), .C2(new_n564), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n628), .A2(new_n627), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT11), .Z(G282));
  INV_X1    g207(.A(new_n631), .ZN(G323));
  NAND2_X1  g208(.A1(new_n494), .A2(new_n464), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n462), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n472), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n463), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT17), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT87), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n661), .A3(new_n665), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n662), .A2(new_n666), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n661), .A2(new_n665), .ZN(new_n672));
  OR3_X1    g247(.A1(new_n671), .A2(new_n664), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n679), .C2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(G160), .A2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(KEYINPUT24), .A2(G34), .ZN(new_n702));
  NOR2_X1   g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT97), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G2084), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT99), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT98), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT26), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n462), .A2(G141), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n472), .A2(G129), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n464), .A2(G105), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n701), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n701), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n708), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n725));
  NAND2_X1  g300(.A1(G103), .A2(G2104), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n462), .A2(G139), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n494), .A2(G127), .ZN(new_n730));
  NAND2_X1  g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n463), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n485), .A2(new_n486), .ZN(new_n735));
  INV_X1    g310(.A(G127), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2105), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n724), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n494), .A2(G139), .A3(new_n463), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n727), .A2(new_n728), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n738), .B2(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n732), .A2(new_n733), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(KEYINPUT96), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n701), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n701), .B2(G33), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(new_n442), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n442), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n723), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT100), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n721), .A2(new_n722), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n701), .A2(G35), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT103), .Z(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n701), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT29), .Z(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G164), .A2(new_n701), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G27), .B2(new_n701), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n760), .B1(new_n443), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n443), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n758), .B2(new_n759), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n767), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n706), .A2(new_n707), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT102), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n701), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n462), .A2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n472), .A2(G128), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(new_n701), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT31), .B(G11), .Z(new_n786));
  INV_X1    g361(.A(G28), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(KEYINPUT30), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT101), .Z(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n642), .B2(new_n701), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n773), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n754), .A2(new_n766), .A3(new_n771), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n767), .A2(G19), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n565), .B2(new_n767), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1341), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n767), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(G299), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n767), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1956), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n794), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n767), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n619), .B2(new_n767), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G1348), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G21), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G168), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1966), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G1348), .B2(new_n805), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n753), .A2(new_n803), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n585), .A2(new_n812), .A3(new_n588), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n585), .B2(new_n588), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G16), .B2(G23), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT33), .B(G1976), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  MUX2_X1   g395(.A(G6), .B(G305), .S(G16), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT32), .B(G1981), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n767), .A2(G22), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT92), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n767), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G1971), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(G1971), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n701), .A2(G25), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n462), .A2(G131), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n472), .A2(G119), .ZN(new_n835));
  OR2_X1    g410(.A1(G95), .A2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n839), .B2(new_n701), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G1986), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n767), .A2(G24), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G290), .B2(G16), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n830), .B2(KEYINPUT34), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT36), .B1(new_n832), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n831), .A4(new_n847), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n811), .B1(new_n849), .B2(new_n852), .ZN(G311));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n852), .ZN(new_n854));
  INV_X1    g429(.A(new_n811), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(G150));
  XOR2_X1   g431(.A(KEYINPUT104), .B(G93), .Z(new_n857));
  NAND3_X1  g432(.A1(new_n553), .A2(new_n501), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n553), .A2(G55), .A3(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n499), .B2(new_n500), .ZN(new_n861));
  AND2_X1   g436(.A1(G80), .A2(G543), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n516), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n858), .A2(new_n859), .A3(new_n866), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n619), .A2(G559), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n561), .A2(new_n563), .A3(new_n864), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n560), .A3(new_n867), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n872), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G860), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n876), .A2(new_n877), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(G145));
  AND3_X1   g457(.A1(new_n740), .A2(new_n783), .A3(new_n746), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n783), .B1(new_n740), .B2(new_n746), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n488), .B1(new_n493), .B2(new_n496), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n493), .A2(new_n496), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n480), .A2(G114), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(G2105), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n472), .A2(G126), .B1(new_n890), .B2(new_n479), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n783), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n734), .A2(new_n739), .A3(new_n724), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT96), .B1(new_n744), .B2(new_n745), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n740), .A2(new_n746), .A3(new_n783), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n718), .B1(new_n886), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n472), .A2(G130), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n463), .A2(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(G142), .B2(new_n462), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n635), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n839), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n885), .B1(new_n883), .B2(new_n884), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n896), .A2(new_n892), .A3(new_n897), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n719), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(KEYINPUT108), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n909), .ZN(new_n913));
  INV_X1    g488(.A(new_n906), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g490(.A(KEYINPUT106), .B(new_n906), .C1(new_n899), .C2(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(G160), .B(new_n642), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n476), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n911), .B(new_n919), .C1(new_n915), .C2(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT107), .B(G37), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT40), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n926));
  INV_X1    g501(.A(new_n924), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n926), .B(new_n927), .C1(new_n921), .C2(new_n922), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(new_n928), .ZN(G395));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n868), .B2(new_n602), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n617), .A2(new_n800), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n617), .A2(new_n800), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n614), .A2(G299), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n617), .A2(new_n800), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n617), .A2(KEYINPUT79), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n615), .B(new_n612), .C1(new_n606), .C2(new_n607), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n625), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n875), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n873), .A2(new_n874), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n619), .A2(new_n625), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n941), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n934), .A2(new_n935), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n946), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT42), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n941), .A2(new_n946), .A3(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n946), .A2(new_n948), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n954), .B(new_n955), .C1(new_n956), .C2(new_n951), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n815), .B1(new_n525), .B2(new_n521), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT73), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(new_n524), .C1(new_n814), .C2(new_n813), .ZN(new_n961));
  XNOR2_X1  g536(.A(G305), .B(G290), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n958), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n953), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G868), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n953), .B2(new_n957), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n931), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n953), .A2(new_n957), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(new_n967), .A3(new_n930), .A4(G868), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n970), .A2(new_n973), .ZN(G295));
  AND2_X1   g549(.A1(new_n970), .A2(new_n973), .ZN(G331));
  AND3_X1   g550(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n976));
  AOI21_X1  g551(.A(G301), .B1(new_n541), .B2(new_n542), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n947), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n535), .A2(new_n536), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT74), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT75), .B1(new_n983), .B2(new_n534), .ZN(new_n984));
  INV_X1    g559(.A(new_n542), .ZN(new_n985));
  OAI21_X1  g560(.A(G171), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n875), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n950), .B1(new_n978), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n947), .B1(new_n976), .B2(new_n977), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n938), .B1(new_n934), .B2(new_n935), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n986), .A2(new_n875), .A3(new_n987), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n937), .A2(new_n939), .A3(new_n933), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n966), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT41), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n932), .B1(new_n937), .B2(new_n939), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n992), .B(new_n990), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n965), .A3(new_n989), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n997), .A3(new_n924), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n989), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n966), .ZN(new_n1004));
  INV_X1    g579(.A(G37), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1002), .B1(new_n1006), .B2(new_n997), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n996), .A2(new_n924), .A3(new_n1001), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1010), .B2(KEYINPUT43), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1004), .A2(new_n997), .A3(new_n1005), .A4(new_n1001), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT111), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1001), .A2(new_n924), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n965), .B1(new_n989), .B2(new_n994), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AND4_X1   g591(.A1(KEYINPUT111), .A2(new_n1016), .A3(KEYINPUT44), .A4(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1013), .B2(new_n1017), .ZN(G397));
  NAND3_X1  g593(.A1(new_n960), .A2(G8), .A3(new_n524), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n960), .A2(KEYINPUT55), .A3(G8), .A4(new_n524), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G164), .B2(G1384), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n887), .B2(new_n891), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT112), .B(G1971), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n892), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1027), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n484), .A2(new_n490), .A3(new_n487), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n490), .B1(new_n484), .B2(new_n487), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n887), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT113), .B(G2090), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1024), .B1(new_n1033), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n813), .A2(new_n814), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT114), .B(G1976), .Z(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n585), .B2(new_n588), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT115), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G288), .A2(KEYINPUT91), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n585), .A2(new_n588), .A3(new_n812), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(G1976), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1050), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n1054), .B2(KEYINPUT52), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n553), .A2(new_n593), .ZN(new_n1067));
  OAI211_X1 g642(.A(G86), .B(new_n501), .C1(new_n507), .C2(new_n508), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n592), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT116), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n594), .A2(new_n595), .A3(new_n1066), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1065), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n594), .A2(new_n595), .A3(new_n1066), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT116), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n592), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT49), .B(new_n1076), .C1(new_n1079), .C2(new_n1066), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1080), .A3(new_n1061), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1051), .A2(new_n1064), .A3(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1076), .B(KEYINPUT117), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G288), .A2(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1046), .A2(new_n1082), .B1(new_n1085), .B2(new_n1050), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1025), .B(G1384), .C1(new_n887), .C2(new_n891), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1025), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1031), .B1(new_n1090), .B2(new_n1027), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1040), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1043), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1027), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1095), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n1043), .A3(new_n1092), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1033), .A2(KEYINPUT118), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(G8), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1023), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1051), .A2(new_n1064), .A3(new_n1081), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1040), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1025), .B1(new_n885), .B2(G1384), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1027), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1966), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1042), .A2(new_n707), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1109), .A2(G286), .A3(new_n1024), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1046), .A3(new_n1104), .A4(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1082), .B1(new_n1023), .B2(new_n1045), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1110), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1086), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1024), .B1(new_n1109), .B2(G168), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1040), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1108), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1089), .A2(KEYINPUT50), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n707), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G286), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1118), .B1(new_n1119), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(G168), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1130), .A2(new_n1118), .A3(G8), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(G8), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT51), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1131), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(G2078), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n489), .A2(new_n491), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1384), .B1(new_n1142), .B2(new_n887), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1125), .B1(new_n1143), .B2(new_n1034), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1139), .A2(new_n1141), .B1(new_n1144), .B2(new_n770), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1026), .A2(new_n443), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1140), .ZN(new_n1147));
  AOI21_X1  g722(.A(G301), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1114), .A2(new_n1103), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1131), .B1(new_n1133), .B2(KEYINPUT51), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1104), .A2(new_n1046), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT45), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1153), .A2(new_n1124), .A3(new_n1088), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1099), .B1(new_n1154), .B2(new_n1031), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1024), .B1(new_n1155), .B2(new_n1087), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1023), .B1(new_n1156), .B2(new_n1100), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1151), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1159));
  NOR2_X1   g734(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1088), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1124), .A2(KEYINPUT123), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n465), .A2(new_n469), .A3(new_n1163), .A4(G40), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n1141), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1144), .A2(new_n770), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1166), .A2(new_n1147), .A3(G301), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1159), .B1(new_n1167), .B2(new_n1148), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(G1956), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT56), .B(G2072), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT57), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n575), .A2(new_n580), .A3(new_n1177), .A4(new_n582), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1175), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(G1348), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1049), .B2(G2067), .ZN(new_n1186));
  INV_X1    g761(.A(G2067), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1028), .A2(new_n1027), .A3(KEYINPUT120), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1183), .B1(new_n944), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .A4(new_n1178), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n1194));
  AND4_X1   g769(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .A4(new_n1178), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1172), .A2(new_n1174), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1183), .A2(new_n1192), .A3(KEYINPUT61), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n616), .A2(new_n1200), .A3(new_n618), .ZN(new_n1201));
  OAI21_X1  g776(.A(KEYINPUT60), .B1(new_n942), .B2(new_n943), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1201), .A2(new_n1202), .A3(new_n1190), .ZN(new_n1203));
  XNOR2_X1  g778(.A(KEYINPUT58), .B(G1341), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1124), .A2(G1996), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1205), .B1(new_n1090), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT59), .B1(new_n1207), .B2(new_n564), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT59), .ZN(new_n1209));
  NOR4_X1   g784(.A1(new_n1153), .A2(G1996), .A3(new_n1088), .A4(new_n1124), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1209), .B(new_n565), .C1(new_n1210), .C2(new_n1205), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  OAI221_X1 g787(.A(KEYINPUT60), .B1(new_n1184), .B2(new_n1189), .C1(new_n942), .C2(new_n943), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1203), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1193), .B1(new_n1199), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT53), .B1(new_n1154), .B2(new_n443), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1218), .B1(new_n1042), .B2(G1961), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1166), .A2(new_n1147), .A3(KEYINPUT125), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1220), .A2(G171), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1144), .A2(new_n770), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1147), .A2(new_n1223), .A3(G301), .A4(new_n1224), .ZN(new_n1225));
  AND2_X1   g800(.A1(new_n1225), .A2(KEYINPUT54), .ZN(new_n1226));
  AOI22_X1  g801(.A1(new_n1168), .A2(new_n1169), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1158), .A2(new_n1170), .A3(new_n1215), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1148), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1152), .A2(new_n1157), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1230), .A2(new_n1231), .A3(new_n1137), .A4(new_n1132), .ZN(new_n1232));
  NAND4_X1  g807(.A1(new_n1117), .A2(new_n1150), .A3(new_n1228), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1160), .A2(new_n1027), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g810(.A(G1996), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n719), .A2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g812(.A(new_n783), .B(G2067), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n718), .A2(G1996), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1240), .ZN(new_n1241));
  OR2_X1    g816(.A1(new_n839), .A2(new_n841), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n839), .A2(new_n841), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(G290), .B(G1986), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1233), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g822(.A1(new_n1234), .A2(G1996), .ZN(new_n1248));
  XNOR2_X1  g823(.A(new_n1248), .B(KEYINPUT46), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1234), .B1(new_n719), .B2(new_n1238), .ZN(new_n1250));
  NOR2_X1   g825(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n1251), .B(KEYINPUT47), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1243), .B1(new_n1240), .B2(new_n1235), .ZN(new_n1253));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1254));
  NOR2_X1   g829(.A1(new_n893), .A2(G2067), .ZN(new_n1255));
  OR3_X1    g830(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1254), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1257));
  AND3_X1   g832(.A1(new_n1256), .A2(new_n1235), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1244), .A2(new_n1235), .ZN(new_n1259));
  NOR3_X1   g834(.A1(new_n1234), .A2(G1986), .A3(G290), .ZN(new_n1260));
  XOR2_X1   g835(.A(new_n1260), .B(KEYINPUT48), .Z(new_n1261));
  AOI211_X1 g836(.A(new_n1252), .B(new_n1258), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1247), .A2(new_n1262), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g838(.A1(new_n923), .A2(new_n924), .ZN(new_n1265));
  INV_X1    g839(.A(G319), .ZN(new_n1266));
  NOR3_X1   g840(.A1(G401), .A2(G227), .A3(new_n1266), .ZN(new_n1267));
  AND3_X1   g841(.A1(new_n697), .A2(new_n698), .A3(new_n1267), .ZN(new_n1268));
  AND3_X1   g842(.A1(new_n1265), .A2(new_n1268), .A3(new_n1007), .ZN(G308));
  NAND3_X1  g843(.A1(new_n1265), .A2(new_n1268), .A3(new_n1007), .ZN(G225));
endmodule


