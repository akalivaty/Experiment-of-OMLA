//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(G50), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n219), .A2(new_n206), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n208), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NOR4_X1   g0024(.A1(new_n217), .A2(new_n218), .A3(new_n221), .A4(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  INV_X1    g0039(.A(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT66), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n220), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n206), .B1(new_n201), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT72), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR3_X1   g0051(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(G33), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n246), .B1(new_n249), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n206), .A3(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n246), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n205), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(new_n247), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT74), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT75), .B1(new_n267), .B2(KEYINPUT9), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n271), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G41), .A2(G45), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(G1), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n280), .A2(new_n281), .A3(G274), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n279), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G222), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G223), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n271), .C1(G77), .C2(new_n294), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n288), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n270), .B(new_n301), .C1(new_n302), .C2(new_n300), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n269), .B2(new_n303), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n266), .C1(G169), .C2(new_n300), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n227), .A2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n294), .B(new_n311), .C1(G226), .C2(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n280), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n275), .A2(G238), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n285), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n322), .A3(G169), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n323), .C1(new_n307), .C2(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n260), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n261), .A2(G68), .A3(new_n262), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n253), .A2(new_n247), .ZN(new_n329));
  INV_X1    g0129(.A(G77), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n256), .A2(new_n330), .B1(new_n206), .B2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n246), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT11), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n327), .B(new_n328), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n333), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n324), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n319), .A2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n336), .B1(new_n319), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n253), .A2(new_n255), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n256), .B1(new_n206), .B2(new_n330), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n246), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n330), .B1(new_n205), .B2(G20), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n261), .A2(new_n348), .B1(new_n330), .B2(new_n260), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n290), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G1698), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G232), .B1(G107), .B2(new_n353), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT73), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n280), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(KEYINPUT73), .A3(new_n356), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n275), .A2(G244), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n285), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n350), .B1(new_n364), .B2(G190), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(G200), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n307), .ZN(new_n368));
  INV_X1    g0168(.A(new_n350), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n338), .A2(new_n343), .A3(new_n367), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n292), .A2(KEYINPUT76), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G33), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT3), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n351), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT76), .B(G33), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n383), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n376), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n353), .B2(new_n206), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n325), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n240), .A2(new_n325), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n253), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n374), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n246), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT3), .ZN(new_n395));
  AOI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n352), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n325), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n293), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT7), .B1(new_n399), .B2(G20), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n394), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n261), .ZN(new_n404));
  INV_X1    g0204(.A(new_n255), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n262), .ZN(new_n406));
  INV_X1    g0206(.A(new_n260), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n404), .A2(new_n406), .B1(new_n407), .B2(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n275), .A2(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n285), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n276), .B2(G1698), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n399), .A2(new_n414), .B1(G33), .B2(G87), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n412), .B(new_n340), .C1(new_n280), .C2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n280), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n302), .B1(new_n417), .B2(new_n411), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND4_X1   g0219(.A1(KEYINPUT78), .A2(new_n403), .A3(new_n409), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n408), .B1(new_n393), .B2(new_n402), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT78), .B1(new_n421), .B2(new_n419), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT17), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n378), .A2(G33), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n292), .A2(KEYINPUT76), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n290), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n291), .B1(new_n427), .B2(KEYINPUT77), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n380), .A2(new_n381), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n375), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n430), .B2(new_n386), .ZN(new_n431));
  INV_X1    g0231(.A(new_n392), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n395), .A2(new_n352), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n397), .A3(new_n206), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G68), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n396), .A2(new_n397), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT16), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n246), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n409), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n412), .B(G179), .C1(new_n280), .C2(new_n415), .ZN(new_n441));
  OAI21_X1  g0241(.A(G169), .B1(new_n417), .B2(new_n411), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n424), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n443), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n419), .B(new_n409), .C1(new_n433), .C2(new_n439), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n423), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n310), .A2(new_n373), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n399), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n383), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n206), .B2(G107), .ZN(new_n457));
  INV_X1    g0257(.A(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT23), .A3(G20), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n455), .A2(new_n206), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n206), .A2(G87), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n353), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n453), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT85), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n453), .A2(new_n460), .A3(new_n467), .A4(new_n463), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n465), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n246), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT86), .B(new_n246), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n246), .B(new_n260), .C1(new_n205), .C2(G33), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n261), .B1(G1), .B2(new_n292), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(G107), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n260), .A2(new_n458), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT25), .Z(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n296), .A2(G250), .ZN(new_n487));
  INV_X1    g0287(.A(G294), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n434), .A2(new_n487), .B1(new_n488), .B2(new_n383), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G257), .A2(G1698), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n434), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n399), .A2(KEYINPUT87), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT88), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n271), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n205), .B(G45), .C1(new_n272), .C2(KEYINPUT5), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n500), .B2(KEYINPUT81), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n271), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n498), .A2(new_n499), .B1(G264), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G274), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n271), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n307), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(G264), .ZN(new_n511));
  INV_X1    g0311(.A(new_n499), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n497), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n370), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n486), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n484), .B1(new_n473), .B2(new_n474), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n302), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G190), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n477), .A2(new_n480), .ZN(new_n522));
  MUX2_X1   g0322(.A(new_n407), .B(new_n522), .S(G97), .Z(new_n523));
  AOI21_X1  g0323(.A(new_n458), .B1(new_n385), .B2(new_n387), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n458), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  XOR2_X1   g0325(.A(G97), .B(G107), .Z(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n330), .B2(new_n253), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n246), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n505), .A2(G257), .B1(new_n508), .B2(new_n504), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n399), .A2(G244), .A3(new_n296), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G244), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n294), .A2(new_n296), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT80), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n354), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n280), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n370), .B1(new_n533), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n538), .A2(new_n537), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(new_n549), .A3(new_n535), .A4(new_n534), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n271), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n532), .A3(new_n307), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n531), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n533), .B2(new_n547), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n532), .A3(G190), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n530), .A4(new_n523), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n407), .A2(G116), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n476), .B2(G116), .ZN(new_n560));
  INV_X1    g0360(.A(G97), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n535), .B(new_n206), .C1(G33), .C2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n246), .C1(new_n206), .C2(G116), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n370), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G270), .B(new_n280), .C1(new_n501), .C2(new_n503), .ZN(new_n567));
  MUX2_X1   g0367(.A(G257), .B(G264), .S(G1698), .Z(new_n568));
  NAND2_X1  g0368(.A1(new_n399), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n353), .A2(G303), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n509), .B(new_n567), .C1(new_n571), .C2(new_n280), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n563), .B(KEYINPUT20), .ZN(new_n574));
  INV_X1    g0374(.A(new_n559), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n478), .B2(new_n454), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n307), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n509), .A2(new_n567), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n280), .B1(new_n569), .B2(new_n570), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n558), .A2(new_n573), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n572), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(new_n577), .C1(new_n340), .C2(new_n572), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n573), .B2(new_n558), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n566), .A2(new_n572), .A3(KEYINPUT84), .A4(KEYINPUT21), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n582), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n399), .A2(new_n206), .A3(G68), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(G87), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n313), .B2(new_n206), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G97), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n592), .A2(new_n593), .B1(new_n256), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n246), .B1(new_n260), .B2(new_n345), .ZN(new_n597));
  INV_X1    g0397(.A(new_n345), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n477), .A2(new_n598), .A3(new_n480), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n599), .A3(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n205), .A2(new_n507), .A3(G45), .ZN(new_n604));
  INV_X1    g0404(.A(G250), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n273), .B2(G1), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n280), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G238), .A2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n540), .B2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n455), .B1(new_n399), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n607), .B1(new_n610), .B2(new_n280), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n307), .B2(new_n611), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n602), .A2(new_n603), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n477), .A2(G87), .A3(new_n480), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(G200), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT83), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n597), .A3(KEYINPUT83), .A4(new_n615), .ZN(new_n620));
  INV_X1    g0420(.A(new_n611), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G190), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n614), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n557), .A2(new_n588), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n452), .A2(new_n521), .A3(new_n625), .ZN(G372));
  NAND3_X1  g0426(.A1(new_n440), .A2(new_n444), .A3(new_n424), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT18), .B1(new_n421), .B2(new_n443), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n338), .B1(new_n342), .B2(new_n372), .ZN(new_n630));
  INV_X1    g0430(.A(new_n450), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT78), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n448), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n421), .A2(KEYINPUT78), .A3(new_n419), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n635), .B2(KEYINPUT17), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n306), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n309), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(KEYINPUT90), .B(new_n309), .C1(new_n637), .C2(new_n638), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n510), .A2(new_n514), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n517), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n557), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n616), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n597), .A2(new_n615), .A3(KEYINPUT89), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n622), .A2(new_n618), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n600), .B2(new_n613), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n646), .A2(new_n520), .A3(new_n647), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT26), .B1(new_n624), .B2(new_n553), .ZN(new_n655));
  INV_X1    g0455(.A(new_n553), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n613), .A2(new_n600), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n452), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n643), .A2(new_n662), .ZN(G369));
  NAND3_X1  g0463(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n644), .A2(new_n577), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n577), .A2(new_n670), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n588), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n516), .B(new_n520), .C1(new_n517), .C2(new_n670), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n516), .B2(new_n670), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n669), .B(KEYINPUT91), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n516), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n644), .A2(new_n669), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n521), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n222), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n590), .A2(new_n591), .A3(new_n454), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n687), .A2(new_n205), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n687), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n689), .A2(KEYINPUT92), .B1(new_n219), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(KEYINPUT92), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT28), .Z(new_n693));
  AOI21_X1  g0493(.A(new_n681), .B1(new_n654), .B2(new_n660), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n651), .A2(new_n652), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n659), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n697), .B2(new_n553), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n659), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n624), .A2(new_n553), .A3(KEYINPUT26), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n669), .B1(new_n654), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n611), .A2(new_n307), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n551), .A2(new_n532), .A3(new_n581), .A4(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n506), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n511), .B1(new_n512), .B2(new_n497), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT30), .B1(new_n711), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n572), .A2(new_n307), .A3(new_n611), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n551), .B2(new_n532), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n513), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n710), .A2(new_n712), .B1(new_n715), .B2(new_n513), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n670), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n516), .A2(new_n625), .A3(new_n520), .A4(new_n680), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n705), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n704), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n693), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n220), .B1(G20), .B2(new_n370), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n686), .A2(new_n353), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n454), .B2(new_n686), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n222), .A2(new_n434), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT93), .Z(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G45), .B2(new_n219), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n243), .A2(G45), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT94), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n259), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n205), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n687), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n340), .A2(new_n302), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n206), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G87), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n206), .A2(new_n307), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n749), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n247), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(G190), .A3(new_n302), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n757), .A2(new_n240), .B1(new_n759), .B2(new_n330), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n340), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n206), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n561), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n302), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n750), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n294), .B1(new_n765), .B2(new_n458), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n756), .A2(new_n760), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n750), .A2(new_n758), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n391), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n754), .A2(KEYINPUT97), .A3(new_n764), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT97), .B1(new_n754), .B2(new_n764), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n767), .B(new_n771), .C1(new_n325), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT98), .Z(new_n776));
  INV_X1    g0576(.A(new_n755), .ZN(new_n777));
  INV_X1    g0577(.A(new_n768), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n777), .A2(G326), .B1(new_n778), .B2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n765), .ZN(new_n781));
  INV_X1    g0581(.A(new_n759), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G311), .A2(new_n782), .B1(new_n752), .B2(G303), .ZN(new_n783));
  INV_X1    g0583(.A(new_n757), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n294), .B1(new_n784), .B2(G322), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(new_n488), .C2(new_n762), .ZN(new_n786));
  INV_X1    g0586(.A(new_n774), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n781), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n776), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n790), .A2(KEYINPUT99), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n732), .B1(new_n790), .B2(KEYINPUT99), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n744), .B(new_n748), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n731), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n673), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT100), .Z(new_n797));
  NOR2_X1   g0597(.A1(new_n673), .A2(G330), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n798), .B(new_n675), .C1(new_n690), .C2(new_n746), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND3_X1  g0601(.A1(new_n368), .A2(new_n371), .A3(new_n670), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n365), .A2(new_n366), .B1(new_n350), .B2(new_n669), .ZN(new_n803));
  INV_X1    g0603(.A(new_n372), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n694), .B(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n748), .B1(new_n807), .B2(new_n725), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n725), .B2(new_n807), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n777), .B1(new_n782), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n811), .B2(new_n757), .C1(new_n774), .C2(new_n254), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(new_n765), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G68), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n247), .B2(new_n751), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT101), .Z(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n399), .B1(new_n820), .B2(new_n768), .C1(new_n240), .C2(new_n762), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n814), .A2(new_n815), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n768), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n765), .A2(new_n591), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(G303), .C2(new_n777), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n787), .A2(G283), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n353), .B1(new_n759), .B2(new_n454), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n757), .A2(new_n488), .B1(new_n751), .B2(new_n458), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n828), .A2(new_n763), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n732), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n748), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n732), .A2(new_n729), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n330), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(new_n806), .C2(new_n730), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n809), .A2(new_n836), .ZN(G384));
  NOR3_X1   g0637(.A1(new_n220), .A2(new_n206), .A3(new_n454), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n527), .B(KEYINPUT102), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT35), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT36), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n219), .A2(new_n330), .A3(new_n389), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n247), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n205), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n667), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n440), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT37), .B1(new_n440), .B2(new_n444), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n852), .A2(new_n633), .A3(new_n634), .A4(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n440), .A2(new_n444), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n850), .A3(new_n448), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n451), .A2(new_n851), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT105), .B1(new_n857), .B2(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n853), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n449), .B1(new_n633), .B2(new_n634), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n860), .A2(new_n629), .A3(new_n631), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n859), .B1(new_n861), .B2(new_n850), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g0666(.A1(new_n633), .A2(new_n852), .A3(new_n634), .A4(new_n850), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n420), .A2(new_n422), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT104), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT16), .B1(new_n870), .B2(KEYINPUT103), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n401), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n439), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n874), .B2(new_n408), .ZN(new_n875));
  INV_X1    g0675(.A(new_n873), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n374), .B1(new_n401), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n402), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n409), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n849), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n444), .A3(new_n879), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n868), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n867), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n636), .B2(new_n447), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT39), .B1(new_n885), .B2(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n866), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n853), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n451), .A2(new_n849), .A3(new_n875), .A4(new_n879), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n883), .A2(new_n884), .A3(new_n864), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT106), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT106), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n324), .A2(new_n337), .A3(new_n670), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n802), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n694), .B2(new_n806), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n337), .A2(new_n669), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n338), .A2(new_n343), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n337), .B(new_n669), .C1(new_n324), .C2(new_n342), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n891), .A2(new_n892), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n909), .A2(new_n910), .B1(new_n629), .B2(new_n667), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n901), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n695), .A2(new_n452), .A3(new_n703), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n643), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n892), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n866), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n723), .A2(new_n721), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n805), .B1(new_n905), .B2(new_n906), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n919), .B(new_n920), .C1(new_n891), .C2(new_n892), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n917), .A2(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n452), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n917), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n452), .A2(new_n919), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n925), .A2(new_n930), .A3(G330), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n915), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n205), .B2(new_n745), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n915), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n848), .B1(new_n933), .B2(new_n934), .ZN(G367));
  INV_X1    g0735(.A(new_n531), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n647), .B1(new_n936), .B2(new_n680), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n553), .B2(new_n680), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n678), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT109), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n521), .A2(new_n938), .A3(new_n683), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n553), .B1(new_n937), .B2(new_n516), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n942), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT108), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n942), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT43), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n653), .B1(new_n651), .B2(new_n670), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n651), .A2(new_n659), .A3(new_n670), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n949), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n941), .A2(new_n957), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n961), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n687), .B(KEYINPUT41), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n684), .A2(new_n938), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT45), .Z(new_n967));
  NAND2_X1  g0767(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n684), .B2(new_n938), .ZN(new_n969));
  NOR2_X1   g0769(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT111), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n969), .A2(new_n972), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n678), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n677), .A2(new_n683), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n521), .A2(new_n683), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n977), .A2(new_n674), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n674), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n967), .A2(new_n679), .A3(new_n973), .A4(new_n974), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n976), .A2(new_n727), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n965), .B1(new_n984), .B2(new_n727), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n962), .B(new_n964), .C1(new_n985), .C2(new_n747), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n738), .A2(new_n233), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n734), .B1(new_n686), .B2(new_n598), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n833), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n732), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n751), .A2(new_n454), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  INV_X1    g0792(.A(new_n762), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(G107), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n787), .A2(G294), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n765), .A2(new_n561), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n759), .A2(new_n780), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G303), .C2(new_n784), .ZN(new_n998));
  INV_X1    g0798(.A(G317), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n755), .A2(new_n823), .B1(new_n768), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n399), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n995), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n816), .A2(G77), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n254), .B2(new_n757), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G143), .B2(new_n777), .ZN(new_n1005));
  INV_X1    g0805(.A(G137), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n751), .A2(new_n240), .B1(new_n768), .B2(new_n1006), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n353), .B(new_n1007), .C1(G50), .C2(new_n782), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n762), .A2(new_n325), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n787), .A2(G159), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1005), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1002), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n989), .B1(new_n990), .B2(new_n1014), .C1(new_n959), .C2(new_n795), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n986), .A2(new_n1015), .ZN(G387));
  OR2_X1    g0816(.A1(new_n677), .A2(new_n795), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n735), .A2(new_n688), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(G107), .B2(new_n222), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n738), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n405), .A2(new_n247), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n273), .B1(new_n325), .B2(new_n330), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n688), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n230), .A2(G45), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n748), .B1(new_n1027), .B2(new_n734), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n787), .A2(new_n405), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n993), .A2(new_n598), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n751), .A2(new_n330), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1031), .A2(new_n996), .A3(new_n434), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n757), .A2(new_n247), .B1(new_n755), .B2(new_n391), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n759), .A2(new_n325), .B1(new_n768), .B2(new_n254), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G116), .A2(new_n816), .B1(new_n778), .B2(G326), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n762), .A2(new_n780), .B1(new_n751), .B2(new_n488), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G322), .A2(new_n777), .B1(new_n782), .B2(G303), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n999), .B2(new_n757), .C1(new_n823), .C2(new_n774), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n434), .B(new_n1037), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1028), .B1(new_n1047), .B2(new_n732), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n982), .A2(new_n747), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n982), .A2(new_n727), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(KEYINPUT112), .A3(new_n687), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n727), .B2(new_n982), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT112), .B1(new_n1050), .B2(new_n687), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(G393));
  NAND3_X1  g0854(.A1(new_n976), .A2(new_n747), .A3(new_n983), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G283), .A2(new_n752), .B1(new_n778), .B2(G322), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n353), .C1(new_n458), .C2(new_n765), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT114), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n757), .A2(new_n823), .B1(new_n755), .B2(new_n999), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n762), .A2(new_n454), .B1(new_n759), .B2(new_n488), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n787), .B2(G303), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n759), .A2(new_n255), .B1(new_n768), .B2(new_n811), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n825), .B(new_n1064), .C1(G68), .C2(new_n752), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n757), .A2(new_n391), .B1(new_n755), .B2(new_n254), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n787), .A2(G50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n434), .B1(new_n993), .B2(G77), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n990), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n738), .A2(new_n237), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n734), .B1(G97), .B2(new_n686), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n833), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1071), .B1(KEYINPUT113), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(KEYINPUT113), .B2(new_n1075), .C1(new_n938), .C2(new_n795), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1055), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT115), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n984), .A2(new_n687), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n976), .A2(new_n983), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1050), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT116), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1084), .A3(new_n1050), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1080), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  AND3_X1   g0888(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n887), .A2(new_n896), .A3(new_n893), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n896), .B1(new_n887), .B2(new_n893), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n694), .A2(new_n806), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n802), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n900), .B1(new_n1093), .B2(new_n907), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n803), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n372), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n902), .B1(new_n702), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n899), .B1(new_n1098), .B2(new_n908), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n917), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1089), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n919), .A2(G330), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n452), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n913), .A2(new_n643), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n724), .A2(new_n806), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(KEYINPUT117), .A3(new_n908), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1089), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n907), .B1(new_n724), .B2(new_n806), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1093), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n806), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n908), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n724), .A2(new_n806), .A3(new_n907), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n1098), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1105), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n899), .B1(new_n903), .B2(new_n908), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n895), .A2(new_n1118), .A3(new_n897), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1102), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1105), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1106), .A2(new_n908), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1089), .B1(new_n1110), .B2(KEYINPUT117), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n903), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1114), .A2(new_n1115), .A3(new_n1098), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1101), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1108), .B1(new_n1119), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1120), .B1(new_n1134), .B2(new_n1118), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1123), .A2(new_n1136), .A3(new_n687), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n747), .B1(new_n1095), .B2(new_n1120), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT118), .B1(new_n1138), .B2(new_n1133), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n746), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT118), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1102), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n833), .B1(new_n255), .B2(new_n834), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n784), .A2(G116), .B1(new_n777), .B2(G283), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n488), .B2(new_n768), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n787), .B2(G107), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n782), .A2(G97), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n753), .A2(new_n1148), .A3(new_n817), .A4(new_n353), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G77), .B2(new_n993), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n294), .B1(new_n768), .B2(new_n1151), .C1(new_n762), .C2(new_n391), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n757), .A2(new_n820), .B1(new_n759), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n755), .A2(new_n1155), .B1(new_n765), .B2(new_n247), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT53), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n751), .B2(new_n254), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n752), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n787), .A2(G137), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1147), .A2(new_n1150), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1144), .B1(new_n990), .B2(new_n1162), .C1(new_n898), .C2(new_n730), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1137), .A2(new_n1143), .A3(new_n1163), .ZN(G378));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n267), .A2(new_n667), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT121), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n310), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n310), .A2(new_n1168), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n928), .B2(new_n705), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n924), .A2(G330), .A3(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1134), .A2(new_n899), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n911), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n901), .A2(new_n911), .A3(new_n1178), .A4(new_n1177), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1176), .A2(new_n729), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n834), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n748), .B1(G50), .B2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT120), .Z(new_n1188));
  OAI22_X1  g0988(.A1(new_n755), .A2(new_n1151), .B1(new_n759), .B2(new_n1006), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n757), .A2(new_n1155), .B1(new_n751), .B2(new_n1153), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G150), .C2(new_n993), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n820), .B2(new_n774), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT119), .Z(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n292), .B(new_n272), .C1(new_n765), .C2(new_n391), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G124), .B2(new_n778), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n434), .A2(new_n272), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1031), .B1(G116), .B2(new_n777), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n784), .A2(G107), .B1(new_n816), .B2(G58), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n598), .A2(new_n782), .B1(new_n778), .B2(G283), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1010), .A4(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1200), .B(new_n1204), .C1(G97), .C2(new_n787), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1200), .B(new_n247), .C1(G33), .C2(G41), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1199), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1188), .B1(new_n1209), .B2(new_n732), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1184), .A2(new_n747), .B1(new_n1185), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1184), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n687), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1184), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT122), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1216), .A2(KEYINPUT122), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n747), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n748), .B1(G68), .B2(new_n1186), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G294), .A2(new_n777), .B1(new_n782), .B2(G107), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n561), .B2(new_n751), .C1(new_n774), .C2(new_n454), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n784), .A2(G283), .B1(new_n778), .B2(G303), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(new_n353), .A3(new_n1003), .A4(new_n1030), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n784), .A2(G137), .B1(new_n777), .B2(G132), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G159), .A2(new_n752), .B1(new_n778), .B2(G128), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n774), .C2(new_n1153), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G150), .A2(new_n782), .B1(new_n816), .B2(G58), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n399), .C1(new_n247), .C2(new_n762), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1225), .A2(new_n1227), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1223), .B1(new_n1233), .B2(new_n732), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n907), .B2(new_n730), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1222), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1221), .A2(new_n1124), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1117), .A2(new_n965), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G381));
  NOR3_X1   g1041(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1087), .A2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1243), .A2(G387), .A3(G381), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT123), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1137), .A2(new_n1143), .A3(new_n1246), .A4(new_n1163), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1244), .B(new_n1248), .C1(new_n1218), .C2(new_n1219), .ZN(G407));
  NAND2_X1  g1049(.A1(new_n668), .A2(G213), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G375), .C2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1253), .B(new_n1254), .ZN(G409));
  INV_X1    g1055(.A(new_n965), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1212), .A2(new_n1256), .A3(new_n1184), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1211), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1245), .A2(new_n1247), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT125), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1211), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1245), .A2(new_n1258), .A3(new_n1262), .A4(new_n1247), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(new_n1237), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n690), .B1(new_n1265), .B2(new_n1237), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1236), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(G384), .B(KEYINPUT126), .Z(new_n1269));
  OR2_X1    g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(KEYINPUT126), .B2(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1264), .A2(new_n1250), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1264), .A2(new_n1250), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1251), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1270), .A2(new_n1271), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1264), .A2(new_n1283), .A3(new_n1250), .A4(new_n1273), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1275), .A2(new_n1281), .A3(new_n1282), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1087), .A2(G387), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n986), .B(new_n1015), .C1(new_n1079), .C2(new_n1086), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(new_n800), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1289), .A3(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1274), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1296), .B(new_n1297), .C1(new_n1295), .C2(new_n1274), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1294), .A2(new_n1298), .ZN(G405));
  OR2_X1    g1099(.A1(new_n1216), .A2(KEYINPUT122), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1217), .A3(new_n1248), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1261), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1292), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1289), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1273), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1291), .A2(new_n1272), .A3(new_n1292), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1302), .B1(new_n1301), .B2(new_n1261), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1304), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1301), .A2(new_n1261), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT127), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1313), .A2(new_n1303), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1311), .A2(new_n1314), .ZN(G402));
endmodule


