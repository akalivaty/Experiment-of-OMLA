//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(KEYINPUT72), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(G902), .C1(new_n189), .C2(new_n190), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT21), .B(G898), .Z(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G122), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT69), .B(G116), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G122), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G128), .B(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT13), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n208), .A2(KEYINPUT13), .A3(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(G134), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT89), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n211), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n205), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n206), .A2(new_n213), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n217), .A2(new_n214), .B1(new_n203), .B2(new_n204), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(G122), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n220));
  INV_X1    g034(.A(new_n201), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n202), .A2(KEYINPUT14), .A3(G122), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(G107), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n218), .A2(new_n224), .A3(KEYINPUT90), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT90), .B1(new_n218), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n216), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT9), .B(G234), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G217), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n229), .A2(new_n230), .A3(G953), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n216), .B(new_n231), .C1(new_n225), .C2(new_n226), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G478), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT15), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(new_n239), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT18), .A2(G131), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n195), .A2(G214), .A3(new_n190), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(G237), .B1(new_n192), .B2(new_n194), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(G143), .A3(G214), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n243), .B1(new_n249), .B2(KEYINPUT86), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n251));
  INV_X1    g065(.A(new_n243), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n246), .A2(new_n251), .A3(new_n252), .A4(new_n248), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G140), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G140), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT85), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n256), .B2(new_n258), .ZN(new_n262));
  OAI21_X1  g076(.A(G146), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n256), .A2(new_n258), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n248), .ZN(new_n269));
  AOI21_X1  g083(.A(G143), .B1(new_n247), .B2(G214), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT17), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n246), .A2(new_n273), .A3(new_n248), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n264), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT16), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n255), .A3(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT76), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n259), .B2(new_n277), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n280), .A3(G146), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G146), .B1(new_n276), .B2(new_n280), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n273), .B1(new_n246), .B2(new_n248), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT17), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n268), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(G113), .B(G122), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(G104), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT88), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  INV_X1    g106(.A(new_n290), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n292), .B(new_n293), .C1(new_n268), .C2(new_n287), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n290), .B(KEYINPUT87), .Z(new_n295));
  AND3_X1   g109(.A1(new_n268), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n291), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G475), .B1(new_n297), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(G475), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT19), .B1(new_n260), .B2(new_n262), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n300), .B(new_n265), .C1(KEYINPUT19), .C2(new_n259), .ZN(new_n301));
  INV_X1    g115(.A(new_n274), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n281), .C1(new_n302), .C2(new_n285), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n293), .B1(new_n268), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n299), .B(new_n236), .C1(new_n296), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT20), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n268), .A2(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n290), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n268), .A2(new_n287), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT20), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n299), .A4(new_n236), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  AND4_X1   g127(.A1(new_n199), .A2(new_n242), .A3(new_n298), .A4(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G210), .B1(G237), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n319));
  XOR2_X1   g133(.A(G110), .B(G122), .Z(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT8), .Z(new_n321));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n322));
  AND2_X1   g136(.A1(KEYINPUT68), .A2(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(KEYINPUT68), .A2(G119), .ZN(new_n324));
  OAI21_X1  g138(.A(G116), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT69), .A2(G116), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT69), .A2(G116), .ZN(new_n327));
  OAI21_X1  g141(.A(G119), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT67), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(KEYINPUT2), .B2(G113), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT2), .A2(G113), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n322), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n332), .A2(new_n334), .B1(KEYINPUT2), .B2(G113), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n325), .A4(new_n328), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n204), .A3(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g158(.A(G101), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n204), .A2(G104), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n348), .A3(new_n204), .A4(G104), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n204), .A2(G104), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n351), .B2(new_n346), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n325), .A2(new_n328), .A3(KEYINPUT5), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(G113), .C1(KEYINPUT5), .C2(new_n325), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n341), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n341), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n321), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G143), .B(G146), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  NOR2_X1   g177(.A1(KEYINPUT0), .A2(G128), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n265), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n245), .A2(G146), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(G128), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT65), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n375), .A3(KEYINPUT1), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(G128), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n368), .A2(new_n369), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n372), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n367), .B1(new_n379), .B2(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n187), .A2(G224), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n359), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n382), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n319), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n341), .A2(new_n354), .A3(new_n356), .ZN(new_n389));
  INV_X1    g203(.A(new_n320), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n338), .A2(new_n340), .B1(new_n337), .B2(new_n329), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n344), .A2(new_n347), .A3(new_n349), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n385), .B(KEYINPUT83), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT84), .A3(new_n383), .A4(new_n359), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n388), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n389), .B1(new_n391), .B2(new_n397), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n320), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n380), .B(new_n381), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n406), .A3(new_n320), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n236), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n318), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n236), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n388), .A2(new_n398), .A3(new_n400), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n317), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n316), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n229), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G469), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n379), .A2(new_n353), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n208), .B1(new_n368), .B2(KEYINPUT1), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n371), .B1(new_n419), .B2(new_n360), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n350), .A3(new_n352), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G137), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G134), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT11), .B1(new_n213), .B2(G137), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT11), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n423), .A3(G134), .ZN(new_n427));
  AOI211_X1 g241(.A(G131), .B(new_n424), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n427), .ZN(new_n429));
  INV_X1    g243(.A(new_n424), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n273), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n422), .A2(KEYINPUT12), .A3(new_n433), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT12), .B1(new_n422), .B2(new_n433), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n435), .B(new_n432), .C1(new_n418), .C2(new_n421), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT82), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n394), .A2(new_n366), .A3(new_n396), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n377), .A2(new_n378), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n371), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n354), .A3(KEYINPUT10), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n421), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n443), .A2(new_n446), .A3(new_n432), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n195), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n439), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n394), .A2(new_n366), .A3(new_n396), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n208), .B1(new_n373), .B2(KEYINPUT65), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n360), .B1(new_n457), .B2(new_n376), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT10), .B1(new_n458), .B2(new_n372), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n448), .B1(new_n459), .B2(new_n353), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n443), .A2(new_n446), .A3(KEYINPUT81), .A4(new_n448), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n433), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n452), .B1(new_n463), .B2(new_n449), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n417), .B(new_n236), .C1(new_n454), .C2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n417), .A2(new_n236), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n449), .B1(new_n440), .B2(new_n441), .ZN(new_n467));
  INV_X1    g281(.A(new_n452), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n463), .A2(new_n453), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(G469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n416), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n314), .A2(new_n414), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n230), .B1(G234), .B2(new_n236), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT24), .B(G110), .ZN(new_n476));
  OAI21_X1  g290(.A(G128), .B1(new_n323), .B2(new_n324), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n208), .A2(G119), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n483));
  OR4_X1    g297(.A1(KEYINPUT23), .A2(new_n323), .A3(new_n324), .A4(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(KEYINPUT23), .A3(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G110), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n476), .C1(new_n480), .C2(new_n481), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n281), .A3(new_n266), .ZN(new_n492));
  OR3_X1    g306(.A1(new_n480), .A2(new_n481), .A3(new_n476), .ZN(new_n493));
  OAI221_X1 g307(.A(new_n493), .B1(new_n487), .B2(new_n486), .C1(new_n283), .C2(new_n282), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT22), .B(G137), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT78), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT25), .B1(new_n505), .B2(new_n236), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n492), .A2(new_n494), .A3(new_n502), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n492), .B2(new_n494), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n500), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n509), .A2(KEYINPUT25), .A3(new_n510), .A4(new_n236), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n475), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n475), .A2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n515), .A2(KEYINPUT79), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(KEYINPUT79), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n366), .B1(new_n428), .B2(new_n431), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n429), .A2(new_n273), .A3(new_n430), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT64), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n423), .B2(G134), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n423), .A2(G134), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n213), .A2(KEYINPUT64), .A3(G137), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n521), .B(KEYINPUT30), .C1(new_n379), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n445), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n521), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n445), .A2(new_n533), .A3(KEYINPUT66), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n379), .B2(new_n529), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n521), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n391), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n247), .A2(G210), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G101), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n391), .A2(new_n534), .A3(new_n521), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT31), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n544), .A2(KEYINPUT31), .A3(new_n548), .A4(new_n549), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n549), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n555), .A2(KEYINPUT28), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n543), .B2(new_n540), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n548), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G472), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n236), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n544), .A2(new_n549), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n560), .C2(new_n559), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n534), .A2(new_n521), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n543), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT74), .A3(new_n549), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n543), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(KEYINPUT28), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n556), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n548), .A2(KEYINPUT29), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n570), .B(new_n236), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n554), .B2(new_n561), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT32), .A3(new_n563), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n566), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n314), .A2(new_n414), .A3(KEYINPUT91), .A4(new_n471), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n474), .A2(new_n520), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AOI22_X1  g400(.A1(new_n552), .A2(new_n553), .B1(new_n560), .B2(new_n559), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n587), .B2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n564), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n519), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n414), .A2(new_n199), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n471), .A3(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n275), .A2(new_n284), .A3(new_n286), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n250), .A2(new_n253), .B1(new_n266), .B2(new_n263), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n290), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n292), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n288), .A2(KEYINPUT88), .A3(new_n290), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n309), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n236), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(G475), .B1(new_n306), .B2(new_n312), .ZN(new_n600));
  AOI21_X1  g414(.A(G478), .B1(new_n235), .B2(new_n236), .ZN(new_n601));
  NOR2_X1   g415(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT92), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n226), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n218), .A2(new_n224), .A3(KEYINPUT90), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n231), .B1(new_n610), .B2(new_n216), .ZN(new_n611));
  INV_X1    g425(.A(new_n234), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n603), .B(new_n607), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n233), .A2(new_n604), .A3(new_n605), .A4(new_n234), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n601), .B1(new_n615), .B2(G478), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n592), .A2(new_n600), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT93), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n242), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n600), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n592), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT35), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  INV_X1    g439(.A(new_n589), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n504), .B1(KEYINPUT36), .B2(new_n499), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n501), .A2(new_n503), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n627), .A2(new_n514), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n513), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n474), .A2(new_n584), .A3(new_n626), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT94), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n487), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  AND2_X1   g450(.A1(new_n583), .A2(new_n471), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n197), .A2(KEYINPUT95), .A3(G900), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT95), .B1(new_n197), .B2(G900), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n191), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n622), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n642), .A2(new_n632), .A3(new_n414), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  AOI21_X1  g459(.A(KEYINPUT32), .B1(new_n581), .B2(new_n563), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n587), .A2(new_n565), .A3(G472), .A4(G902), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n567), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n560), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n573), .A2(new_n575), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n236), .B1(new_n651), .B2(new_n548), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT96), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT25), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n515), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n511), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n630), .B1(new_n659), .B2(new_n475), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n600), .A2(new_n242), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n315), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n640), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n471), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT40), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n410), .A2(new_n413), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n656), .A2(new_n663), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  AOI211_X1 g485(.A(new_n602), .B(new_n606), .C1(new_n233), .C2(new_n234), .ZN(new_n672));
  INV_X1    g486(.A(new_n614), .ZN(new_n673));
  OAI211_X1 g487(.A(G478), .B(new_n236), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n601), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n298), .A2(new_n313), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n414), .A2(new_n676), .A3(new_n640), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n660), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n600), .A2(new_n616), .A3(new_n641), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT99), .A3(new_n414), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n679), .A2(new_n583), .A3(new_n471), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  AOI21_X1  g497(.A(new_n519), .B1(new_n648), .B2(new_n580), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n236), .B1(new_n454), .B2(new_n464), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n415), .A3(new_n465), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n415), .A4(new_n465), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n199), .A2(new_n689), .A3(new_n414), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n684), .A2(new_n676), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  INV_X1    g508(.A(new_n622), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n520), .A3(new_n583), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NOR3_X1   g511(.A1(new_n401), .A2(new_n318), .A3(new_n409), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n317), .B1(new_n411), .B2(new_n412), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n315), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n660), .A2(new_n700), .A3(new_n687), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n583), .A3(new_n314), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND2_X1  g517(.A1(new_n577), .A2(new_n560), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n554), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n563), .A4(new_n236), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n552), .A2(new_n553), .B1(new_n560), .B2(new_n577), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n563), .A2(new_n236), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT101), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n588), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n519), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n691), .A2(new_n712), .A3(new_n661), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NAND2_X1  g528(.A1(new_n676), .A2(new_n640), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n680), .A2(new_n588), .A3(new_n707), .A4(new_n710), .ZN(new_n719));
  INV_X1    g533(.A(new_n687), .ZN(new_n720));
  INV_X1    g534(.A(new_n475), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n658), .B2(new_n511), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n720), .B(new_n414), .C1(new_n722), .C2(new_n630), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n718), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NAND4_X1  g540(.A1(new_n410), .A2(new_n413), .A3(new_n415), .A4(new_n315), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n465), .B2(new_n470), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n465), .A2(KEYINPUT103), .A3(new_n470), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n465), .A2(KEYINPUT103), .A3(new_n470), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n730), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT104), .B1(new_n736), .B2(new_n727), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n684), .A3(new_n680), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n715), .B1(new_n734), .B2(new_n737), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n566), .A2(new_n743), .A3(new_n582), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT106), .B1(new_n646), .B2(new_n647), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n580), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n520), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NAND3_X1  g563(.A1(new_n738), .A2(new_n684), .A3(new_n642), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND3_X1  g565(.A1(new_n410), .A2(new_n315), .A3(new_n413), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n626), .A2(new_n660), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n298), .A2(new_n313), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n754), .B2(new_n616), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n754), .A2(KEYINPUT43), .A3(new_n616), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n469), .B(KEYINPUT45), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  INV_X1    g575(.A(new_n466), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n764), .B(G469), .C1(new_n760), .C2(G902), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n465), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n415), .ZN(new_n767));
  INV_X1    g581(.A(new_n665), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT107), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n755), .A4(new_n756), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n766), .A2(new_n771), .A3(new_n415), .A4(new_n665), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n759), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n767), .B(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n752), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n520), .A2(new_n583), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n715), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n255), .ZN(G42));
  NAND2_X1  g595(.A1(new_n686), .A2(new_n465), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n754), .A3(new_n616), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g599(.A(new_n782), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n316), .A3(new_n669), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n655), .A3(new_n520), .A4(new_n415), .ZN(new_n789));
  INV_X1    g603(.A(new_n191), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n756), .A2(new_n790), .A3(new_n755), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n728), .A2(new_n786), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n520), .A3(new_n746), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT48), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT117), .Z(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(KEYINPUT48), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT116), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n188), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n767), .B(KEYINPUT47), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n416), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n752), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n791), .A2(new_n519), .A3(new_n711), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n792), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n519), .A2(new_n191), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n655), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n655), .A2(KEYINPUT113), .A3(new_n808), .A4(new_n809), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n600), .A3(new_n616), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n711), .A2(new_n660), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n793), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n806), .A2(new_n720), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n669), .A2(new_n315), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(KEYINPUT50), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n806), .A2(new_n720), .A3(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n807), .A2(new_n814), .A3(new_n816), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n799), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n817), .A2(new_n414), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n416), .B1(new_n648), .B2(new_n653), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n414), .A2(new_n661), .A3(new_n640), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n660), .A3(new_n733), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n725), .A2(new_n831), .A3(new_n644), .A4(new_n682), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n717), .A2(new_n724), .B1(new_n637), .B2(new_n643), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n682), .A4(new_n831), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n692), .A2(new_n696), .A3(new_n702), .A4(new_n713), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n748), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n676), .A2(KEYINPUT108), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT108), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n600), .B2(new_n616), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n622), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n590), .A2(new_n844), .A3(new_n471), .A4(new_n591), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n585), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n754), .A2(new_n621), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n752), .A2(new_n641), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n583), .A2(new_n471), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n719), .B1(new_n734), .B2(new_n737), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n632), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n846), .A2(new_n852), .A3(new_n633), .A4(new_n750), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n840), .A2(new_n853), .A3(KEYINPUT109), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n692), .A2(new_n696), .A3(new_n702), .A4(new_n713), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n747), .B2(new_n741), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n750), .A2(new_n585), .A3(new_n633), .A4(new_n845), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n738), .A2(new_n716), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n660), .B1(new_n859), .B2(new_n849), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n855), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n838), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT53), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT109), .B1(new_n840), .B2(new_n853), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n855), .A3(new_n861), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n836), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n837), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n840), .A2(new_n853), .A3(new_n868), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n871), .A3(new_n869), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n837), .B1(new_n865), .B2(new_n866), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n875), .B(new_n876), .C1(new_n877), .C2(KEYINPUT53), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n827), .A2(new_n828), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n814), .A2(new_n816), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT112), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n819), .B2(new_n822), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n823), .A2(KEYINPUT112), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n880), .B(KEYINPUT114), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n814), .A2(new_n816), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n805), .A2(new_n806), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(new_n800), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n812), .A2(new_n676), .A3(new_n813), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n879), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n789), .B1(new_n893), .B2(new_n894), .ZN(G75));
  NAND2_X1  g709(.A1(new_n404), .A2(new_n407), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT118), .Z(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  OAI21_X1  g712(.A(new_n875), .B1(new_n877), .B2(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G210), .A3(G902), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  INV_X1    g715(.A(new_n405), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n405), .ZN(new_n907));
  INV_X1    g721(.A(new_n898), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n195), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n905), .A2(new_n910), .A3(new_n912), .ZN(G51));
  NAND2_X1  g727(.A1(new_n762), .A2(KEYINPUT57), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n762), .A2(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n878), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n914), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n464), .B2(new_n454), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n899), .A2(G469), .A3(G902), .A4(new_n760), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT119), .Z(new_n922));
  AOI21_X1  g736(.A(new_n911), .B1(new_n920), .B2(new_n922), .ZN(G54));
  NAND4_X1  g737(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n924));
  INV_X1    g738(.A(new_n310), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n911), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n873), .B2(new_n878), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n672), .A2(new_n673), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n912), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n932), .B(new_n930), .C1(new_n916), .C2(new_n878), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT120), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n868), .B1(new_n854), .B2(new_n862), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n871), .A2(new_n869), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n937), .A2(new_n938), .B1(new_n877), .B2(new_n868), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n878), .B1(new_n939), .B2(new_n876), .ZN(new_n940));
  INV_X1    g754(.A(new_n930), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n932), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n933), .B(new_n941), .C1(new_n917), .C2(new_n918), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(new_n944), .A3(new_n912), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n936), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT60), .Z(new_n949));
  AND2_X1   g763(.A1(new_n899), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n629), .A3(new_n627), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n516), .A2(new_n517), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n951), .B(new_n912), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n950), .A2(new_n953), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(KEYINPUT61), .A3(new_n912), .A4(new_n951), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(G66));
  AOI21_X1  g773(.A(new_n187), .B1(new_n198), .B2(G224), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n839), .A2(new_n633), .A3(new_n846), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n195), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n897), .B1(G898), .B2(new_n195), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  NAND2_X1  g779(.A1(new_n536), .A2(new_n542), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n300), .B1(KEYINPUT19), .B2(new_n259), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n196), .A2(G900), .ZN(new_n969));
  INV_X1    g783(.A(new_n780), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n769), .A2(new_n414), .A3(new_n661), .A4(new_n772), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n746), .A2(new_n520), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n750), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n773), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n834), .A2(new_n682), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n970), .A2(new_n975), .A3(new_n748), .A4(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n968), .B(new_n969), .C1(new_n978), .C2(new_n196), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n670), .A2(new_n977), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n670), .A2(new_n977), .A3(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n666), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n684), .A2(new_n985), .A3(new_n777), .A4(new_n844), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n773), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT123), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n773), .A2(new_n989), .A3(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n780), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n196), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n979), .B1(new_n968), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n992), .ZN(new_n996));
  INV_X1    g810(.A(new_n968), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(KEYINPUT124), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n992), .B2(new_n968), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n994), .B(KEYINPUT125), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n979), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  NAND2_X1  g822(.A1(new_n984), .A2(new_n991), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n961), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n650), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n978), .B2(new_n961), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n560), .A3(new_n649), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n912), .A3(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n568), .B(KEYINPUT127), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n939), .B1(new_n550), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1008), .B2(new_n1016), .ZN(G57));
endmodule


