//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n464), .B2(G101), .ZN(new_n465));
  AND4_X1   g040(.A1(KEYINPUT67), .A2(new_n459), .A3(G101), .A4(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT68), .Z(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G136), .A3(new_n459), .ZN(new_n474));
  INV_X1    g049(.A(G100), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n475), .A2(new_n459), .A3(KEYINPUT69), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n475), .B2(new_n459), .ZN(new_n477));
  OAI221_X1 g052(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n459), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n474), .A2(new_n478), .A3(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT70), .A2(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n459), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n473), .A2(new_n494), .A3(G138), .A4(new_n459), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n497), .A3(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n506), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AND2_X1   g091(.A1(new_n503), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n511), .A2(G543), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G52), .Z(new_n532));
  OAI22_X1  g107(.A1(new_n512), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n529), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  XOR2_X1   g110(.A(KEYINPUT74), .B(G43), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n509), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n512), .B2(new_n538), .C1(new_n539), .C2(new_n505), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT75), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n517), .A2(G81), .B1(new_n509), .B2(new_n536), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n542), .B(new_n543), .C1(new_n505), .C2(new_n539), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n509), .A2(new_n552), .A3(G53), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n509), .B2(G53), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n512), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(KEYINPUT76), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n505), .B1(new_n558), .B2(KEYINPUT76), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  NAND2_X1  g139(.A1(new_n509), .A2(G49), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n503), .ZN(new_n568));
  INV_X1    g143(.A(G74), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n505), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n505), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n509), .A2(G48), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  XOR2_X1   g154(.A(KEYINPUT77), .B(G85), .Z(new_n580));
  AOI22_X1  g155(.A1(new_n517), .A2(new_n580), .B1(G47), .B2(new_n509), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n505), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(new_n517), .A2(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n568), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n591), .A2(new_n592), .B1(new_n593), .B2(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(KEYINPUT78), .B2(new_n593), .ZN(G284));
  XOR2_X1   g170(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n592), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G168), .B2(new_n592), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G168), .B2(new_n592), .ZN(G280));
  INV_X1    g174(.A(new_n591), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n545), .A2(new_n592), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT11), .Z(G282));
  INV_X1    g181(.A(new_n605), .ZN(G323));
  NAND2_X1  g182(.A1(new_n473), .A2(new_n459), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n463), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(KEYINPUT13), .B1(KEYINPUT80), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT13), .B2(new_n611), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n614), .A2(KEYINPUT80), .A3(new_n612), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(KEYINPUT80), .B2(new_n612), .ZN(new_n616));
  MUX2_X1   g191(.A(G99), .B(G111), .S(G2105), .Z(new_n617));
  AOI22_X1  g192(.A1(new_n481), .A2(G123), .B1(new_n617), .B2(G2104), .ZN(new_n618));
  INV_X1    g193(.A(G135), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n608), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n615), .A2(new_n616), .A3(new_n621), .ZN(G156));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2427), .ZN(new_n626));
  INV_X1    g201(.A(G2430), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n642), .B(KEYINPUT17), .Z(new_n646));
  INV_X1    g221(.A(new_n641), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  INV_X1    g224(.A(new_n640), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n641), .B2(new_n642), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n645), .B(new_n648), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n663), .A2(new_n664), .A3(new_n660), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n663), .B1(new_n664), .B2(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n669), .B(new_n671), .Z(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  NOR2_X1   g252(.A1(G16), .A2(G23), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n571), .B(KEYINPUT87), .Z(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  NOR2_X1   g257(.A1(G6), .A2(G16), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n578), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  NOR2_X1   g262(.A1(G16), .A2(G22), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G166), .B2(G16), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT88), .B(G1971), .Z(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  NOR3_X1   g266(.A1(new_n682), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n696));
  OR2_X1    g271(.A1(G16), .A2(G24), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(G290), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT84), .B(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  MUX2_X1   g278(.A(G95), .B(G107), .S(G2105), .Z(new_n704));
  AOI22_X1  g279(.A1(new_n481), .A2(G119), .B1(new_n704), .B2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(G131), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n608), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT85), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  AOI211_X1 g287(.A(new_n701), .B(new_n712), .C1(new_n700), .C2(new_n699), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n694), .A2(new_n695), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n702), .A2(G35), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n702), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G2090), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(G2090), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NAND2_X1  g300(.A1(G160), .A2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT24), .B(G34), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n702), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G168), .B2(G16), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1966), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n698), .A2(G19), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n545), .B2(new_n698), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G1341), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n731), .A2(new_n735), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n698), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G1341), .B2(new_n738), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n460), .A2(new_n461), .ZN(new_n747));
  INV_X1    g322(.A(G127), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n464), .A2(G103), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT25), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n464), .A2(new_n755), .A3(G103), .ZN(new_n756));
  INV_X1    g331(.A(G139), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n756), .C1(new_n608), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT90), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(KEYINPUT90), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n752), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G33), .B(new_n761), .S(G29), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  NOR2_X1   g339(.A1(G4), .A2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n600), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT30), .B(G28), .Z(new_n771));
  OAI221_X1 g346(.A(new_n770), .B1(G29), .B2(new_n771), .C1(new_n620), .C2(new_n702), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n481), .A2(G129), .ZN(new_n773));
  INV_X1    g348(.A(G141), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n608), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G105), .B2(new_n464), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G32), .B(new_n781), .S(G29), .Z(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  AOI21_X1  g358(.A(new_n772), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n784), .B1(new_n782), .B2(new_n783), .C1(new_n730), .C2(new_n725), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n698), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n698), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n733), .A2(G1966), .ZN(new_n790));
  MUX2_X1   g365(.A(G104), .B(G116), .S(G2105), .Z(new_n791));
  AOI22_X1  g366(.A1(new_n481), .A2(G128), .B1(new_n791), .B2(G2104), .ZN(new_n792));
  INV_X1    g367(.A(G140), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n608), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n702), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G2067), .Z(new_n799));
  INV_X1    g374(.A(new_n702), .ZN(new_n800));
  NAND2_X1  g375(.A1(G164), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G27), .B2(new_n800), .ZN(new_n802));
  INV_X1    g377(.A(G2078), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n799), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G1348), .B2(new_n766), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n768), .A2(new_n789), .A3(new_n790), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n740), .A2(new_n745), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n716), .A2(new_n717), .A3(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n600), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n509), .A2(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n512), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n505), .B1(new_n818), .B2(KEYINPUT97), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n545), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n540), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n813), .B(new_n826), .Z(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n823), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n761), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n781), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n493), .A2(new_n495), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n484), .B(KEYINPUT98), .C1(new_n489), .C2(new_n490), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n488), .ZN(new_n840));
  NOR2_X1   g415(.A1(KEYINPUT70), .A2(G114), .ZN(new_n841));
  OAI21_X1  g416(.A(G2105), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n490), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT98), .B1(new_n844), .B2(new_n484), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT99), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n491), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n837), .A4(new_n838), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n794), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n836), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n610), .B(new_n707), .Z(new_n854));
  MUX2_X1   g429(.A(G106), .B(G118), .S(G2105), .Z(new_n855));
  AOI22_X1  g430(.A1(new_n481), .A2(G130), .B1(new_n855), .B2(G2104), .ZN(new_n856));
  INV_X1    g431(.A(G142), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n608), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n854), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n836), .A2(new_n852), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n853), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n853), .A2(new_n863), .A3(new_n859), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n853), .A2(new_n860), .ZN(new_n865));
  INV_X1    g440(.A(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G160), .B(G162), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n620), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n861), .A2(new_n870), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n873), .B2(new_n867), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT102), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n877), .A2(KEYINPUT40), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT40), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(G395));
  NOR2_X1   g456(.A1(new_n823), .A2(G868), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n600), .A2(new_n601), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n826), .B(new_n883), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n600), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n591), .A2(new_n562), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n891), .B2(KEYINPUT41), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n884), .A2(new_n887), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT42), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G290), .B(KEYINPUT104), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(new_n679), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n679), .ZN(new_n902));
  XNOR2_X1  g477(.A(G303), .B(new_n578), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n899), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n882), .B1(new_n908), .B2(G868), .ZN(G295));
  AOI21_X1  g484(.A(new_n882), .B1(new_n908), .B2(G868), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  XNOR2_X1  g486(.A(G168), .B(G301), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(new_n826), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n826), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n886), .A3(new_n885), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n905), .A2(new_n919), .A3(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n913), .A2(new_n887), .A3(new_n914), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n913), .A2(new_n914), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n907), .B(new_n924), .C1(new_n925), .C2(new_n892), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n925), .A2(new_n892), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT105), .B1(new_n932), .B2(new_n924), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT105), .B(new_n924), .C1(new_n925), .C2(new_n892), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n921), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n930), .B(new_n931), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n911), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n923), .B2(new_n928), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n930), .B(KEYINPUT43), .C1(new_n933), .C2(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(G397));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n846), .A2(new_n942), .A3(new_n850), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT107), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n467), .A2(new_n470), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n944), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n781), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT108), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n781), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n949), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n794), .B(G2067), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n948), .A2(KEYINPUT109), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT109), .B1(new_n948), .B2(new_n955), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n707), .B(new_n711), .Z(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n948), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n952), .A2(new_n958), .A3(new_n960), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n948), .A2(new_n955), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n953), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n950), .B(KEYINPUT46), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n944), .A2(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n946), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n709), .A2(new_n711), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT125), .Z(new_n976));
  NAND3_X1  g551(.A1(new_n952), .A2(new_n958), .A3(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n794), .A2(G2067), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(G305), .A2(G1981), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT114), .B(G86), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n575), .B1(new_n512), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(G1981), .B1(new_n574), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT49), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n946), .B(new_n942), .C1(new_n839), .C2(new_n845), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(KEYINPUT49), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n679), .A2(G1976), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT52), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n571), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n992), .B2(new_n994), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n990), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n942), .A4(new_n850), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n481), .A2(G126), .B1(new_n842), .B2(new_n843), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n837), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n942), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n947), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1971), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n848), .A2(new_n837), .A3(new_n838), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT50), .B1(new_n1007), .B2(new_n942), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n946), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n1006), .A2(KEYINPUT110), .B1(G2090), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(KEYINPUT111), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1014), .B2(KEYINPUT111), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n1018));
  OAI211_X1 g593(.A(G303), .B(G8), .C1(new_n1018), .C2(KEYINPUT55), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(KEYINPUT55), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1019), .B(new_n1020), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT117), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1015), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1004), .B(new_n942), .C1(new_n839), .C2(new_n845), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT45), .B1(G164), .B2(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1966), .B1(new_n1026), .B2(new_n946), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n942), .B1(new_n839), .B2(new_n845), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n947), .B1(new_n1030), .B2(new_n1009), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1027), .A2(KEYINPUT116), .B1(new_n1031), .B2(new_n725), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n947), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(G1966), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1016), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n999), .A2(new_n1023), .A3(G168), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1022), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT63), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(new_n1021), .ZN(new_n1041));
  INV_X1    g616(.A(new_n990), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G288), .A2(G1976), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT115), .Z(new_n1044));
  OAI21_X1  g619(.A(new_n981), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1041), .A2(new_n999), .B1(new_n988), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(G2078), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1034), .A2(KEYINPUT53), .A3(new_n803), .ZN(new_n1051));
  INV_X1    g626(.A(G1961), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1011), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G168), .A2(new_n1016), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(KEYINPUT51), .C1(new_n1036), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1026), .A2(new_n946), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n725), .B(new_n946), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1035), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT51), .B(G8), .C1(new_n1067), .C2(G286), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1070), .B(new_n1071), .C1(new_n1016), .C2(G168), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1036), .A2(G286), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(KEYINPUT62), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT62), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1059), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n1054), .B2(G171), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1000), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n946), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n973), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1082), .B2(G171), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1057), .B(new_n1058), .C1(G171), .C2(new_n1082), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1000), .A2(new_n1005), .A3(new_n949), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n987), .A2(KEYINPUT119), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1007), .A2(new_n1089), .A3(new_n942), .A4(new_n946), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT58), .B(G1341), .Z(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n545), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT121), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(new_n545), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(KEYINPUT59), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1093), .B2(new_n545), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n541), .A2(new_n544), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT121), .B(new_n1101), .C1(new_n1087), .C2(new_n1092), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT56), .B(G2072), .Z(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1000), .A2(new_n1005), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1003), .A2(new_n1029), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1007), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1956), .B1(new_n1111), .B2(new_n946), .ZN(new_n1112));
  INV_X1    g687(.A(new_n555), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1113), .A2(new_n553), .B1(new_n517), .B2(G91), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n558), .A2(KEYINPUT76), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G651), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1115), .C1(new_n1117), .C2(new_n559), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT57), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n562), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1108), .A2(new_n1112), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1121), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1111), .A2(new_n946), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1123), .B1(new_n1126), .B2(new_n1107), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1104), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1121), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1123), .A3(new_n1107), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT61), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1098), .A2(new_n1103), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(G2067), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1133), .A2(KEYINPUT120), .B1(new_n1011), .B2(new_n764), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1140), .B(G2067), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1031), .A2(G1348), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n591), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT60), .A4(new_n591), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT122), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n600), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1132), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1136), .A2(new_n600), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1122), .B1(new_n1151), .B2(new_n1129), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1078), .B(new_n1086), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1153));
  OR3_X1    g728(.A1(new_n1070), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1077), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1124), .A2(G2090), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1156), .B2(new_n1006), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n998), .B(new_n1041), .C1(new_n1021), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1047), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n948), .B1(new_n961), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n952), .A2(new_n1161), .A3(new_n958), .A4(new_n960), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n980), .B1(new_n1159), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g738(.A1(new_n877), .A2(new_n878), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n654), .A2(G319), .ZN(new_n1166));
  OAI211_X1 g740(.A(new_n676), .B(new_n638), .C1(KEYINPUT127), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g741(.A(new_n1167), .B1(KEYINPUT127), .B2(new_n1166), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n938), .A3(new_n939), .A4(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


