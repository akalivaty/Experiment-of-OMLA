//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n476));
  INV_X1    g051(.A(G100), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n463), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n483), .B2(G138), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n465), .A2(new_n467), .A3(new_n487), .A4(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n463), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(G164));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n504), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n501), .A2(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n499), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  INV_X1    g088(.A(new_n501), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G51), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n505), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n504), .A2(new_n506), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(KEYINPUT72), .B(new_n527), .C1(new_n509), .C2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n496), .A2(new_n500), .A3(G89), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT72), .B1(new_n531), .B2(new_n527), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n515), .B(new_n522), .C1(new_n530), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n501), .A2(new_n535), .B1(new_n509), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n498), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n518), .B2(new_n520), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n504), .A2(new_n506), .A3(new_n519), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n519), .B1(new_n504), .B2(new_n506), .ZN(new_n549));
  OAI21_X1  g124(.A(G56), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(KEYINPUT73), .A3(new_n545), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(G651), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n501), .A2(new_n553), .B1(new_n509), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  XOR2_X1   g136(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G188));
  XNOR2_X1  g140(.A(new_n509), .B(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n496), .A2(G65), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n498), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n501), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n500), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n567), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n566), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n514), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(new_n496), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n514), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n589));
  AOI211_X1 g164(.A(KEYINPUT77), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n566), .B2(G86), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n586), .B1(new_n590), .B2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n498), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n501), .A2(new_n596), .B1(new_n509), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n566), .A2(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n583), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n514), .B2(G54), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n566), .A2(new_n608), .A3(G92), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT78), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G91), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n588), .B2(new_n589), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n574), .A2(new_n575), .ZN(new_n617));
  NOR3_X1   g192(.A1(new_n616), .A2(new_n617), .A3(new_n570), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n614), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n614), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n611), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n610), .B(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(G868), .B1(new_n624), .B2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n483), .A2(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n481), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n483), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2451), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  AOI21_X1  g235(.A(KEYINPUT18), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  MUX2_X1   g236(.A(new_n658), .B(new_n653), .S(new_n661), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n678), .C1(new_n676), .C2(new_n675), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT82), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT22), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G35), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G162), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G2090), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT93), .ZN(new_n692));
  INV_X1    g267(.A(G1961), .ZN(new_n693));
  NAND2_X1  g268(.A1(G171), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G5), .B2(G16), .ZN(new_n695));
  OAI22_X1  g270(.A1(new_n690), .A2(G2090), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  OR2_X1    g272(.A1(KEYINPUT24), .A2(G34), .ZN(new_n698));
  NAND2_X1  g273(.A1(KEYINPUT24), .A2(G34), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n687), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G160), .B2(new_n687), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT90), .Z(new_n702));
  AOI21_X1  g277(.A(new_n696), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G4), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n611), .B2(G16), .ZN(new_n705));
  INV_X1    g280(.A(G1348), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G21), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G168), .B2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT91), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G1966), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n692), .A2(new_n703), .A3(new_n707), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n483), .A2(G139), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n463), .ZN(new_n718));
  MUX2_X1   g293(.A(G33), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2072), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT31), .B(G11), .Z(new_n721));
  INV_X1    g296(.A(new_n702), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G2084), .ZN(new_n723));
  NAND2_X1  g298(.A1(G164), .A2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G27), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2078), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(G128), .A2(new_n481), .B1(new_n483), .B2(G140), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n729));
  NOR2_X1   g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT88), .Z(new_n731));
  OAI21_X1  g306(.A(new_n728), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n687), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(G29), .A2(G32), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n481), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n468), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n743), .C1(new_n744), .C2(G2105), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n687), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n695), .A2(new_n693), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n723), .A2(new_n727), .A3(new_n739), .A4(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT94), .B(KEYINPUT23), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n708), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n618), .B2(new_n708), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(G28), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT30), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n725), .A2(new_n726), .B1(new_n687), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n759), .B1(new_n687), .B2(new_n636), .C1(new_n746), .C2(new_n747), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n713), .A2(new_n720), .A3(new_n749), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n708), .A2(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n558), .B2(new_n708), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT87), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT86), .B(G1341), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n761), .B(new_n766), .C1(G1966), .C2(new_n711), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  MUX2_X1   g343(.A(G6), .B(G305), .S(G16), .Z(new_n769));
  XOR2_X1   g344(.A(KEYINPUT32), .B(G1981), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n708), .A2(G22), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n708), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1971), .Z(new_n774));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G16), .B2(G23), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n775), .A2(G16), .A3(G23), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n776), .B(new_n777), .C1(G288), .C2(new_n708), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n771), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G24), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n599), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT83), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G1986), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(G1986), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT35), .B(G1991), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n481), .A2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n483), .A2(G131), .ZN(new_n791));
  NOR2_X1   g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G25), .B(new_n794), .S(G29), .Z(new_n795));
  AOI211_X1 g370(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n783), .B(new_n796), .C1(new_n789), .C2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT36), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n768), .A2(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  NAND2_X1  g375(.A1(G80), .A2(G543), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n521), .B2(G67), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT98), .B1(new_n803), .B2(new_n498), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  INV_X1    g380(.A(G93), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n501), .A2(new_n805), .B1(new_n509), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(G67), .B1(new_n548), .B2(new_n549), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(new_n801), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n810), .A2(new_n811), .A3(G651), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n804), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n611), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT39), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n811), .B1(new_n810), .B2(G651), .ZN(new_n818));
  AOI211_X1 g393(.A(KEYINPUT98), .B(new_n498), .C1(new_n809), .C2(new_n801), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n557), .A2(new_n820), .A3(new_n808), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n813), .A2(new_n556), .A3(new_n552), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n817), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n815), .B1(new_n827), .B2(G860), .ZN(G145));
  XNOR2_X1  g403(.A(G160), .B(new_n636), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n485), .ZN(new_n830));
  XNOR2_X1  g405(.A(G164), .B(new_n718), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n794), .B(new_n745), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n483), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n481), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n463), .A2(G118), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n834), .B(new_n835), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n832), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n629), .B(new_n732), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n843), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g423(.A(G288), .B(G303), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G290), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(G305), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n624), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n823), .Z(new_n854));
  AND2_X1   g429(.A1(new_n603), .A2(new_n609), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n855), .A2(KEYINPUT100), .A3(new_n618), .A4(new_n607), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g432(.A1(G299), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n618), .A2(KEYINPUT100), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n859), .A3(new_n610), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT41), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n853), .B(new_n823), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n868), .B1(new_n867), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n852), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n867), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n851), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n878), .A3(G868), .ZN(new_n879));
  INV_X1    g454(.A(new_n813), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT101), .B1(new_n880), .B2(G868), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n882), .B(new_n886), .C1(new_n883), .C2(new_n879), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G295));
  NAND2_X1  g463(.A1(new_n884), .A2(KEYINPUT103), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n882), .B(new_n890), .C1(new_n883), .C2(new_n879), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n893));
  XNOR2_X1  g468(.A(G301), .B(G286), .ZN(new_n894));
  AND4_X1   g469(.A1(KEYINPUT104), .A2(new_n894), .A3(new_n821), .A4(new_n822), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n894), .A2(new_n821), .A3(new_n822), .ZN(new_n896));
  NAND2_X1  g471(.A1(G168), .A2(G301), .ZN(new_n897));
  NAND2_X1  g472(.A1(G171), .A2(G286), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n821), .A2(new_n822), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n896), .A2(new_n899), .A3(KEYINPUT104), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n865), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n896), .A2(new_n899), .A3(KEYINPUT105), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n899), .B2(KEYINPUT105), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n861), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n905), .B2(new_n852), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n870), .B1(new_n900), .B2(new_n895), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n862), .A2(new_n909), .A3(new_n864), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n861), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(new_n910), .A3(new_n903), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(new_n870), .C1(new_n900), .C2(new_n895), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n915), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT108), .B1(new_n915), .B2(new_n851), .ZN(new_n917));
  OAI211_X1 g492(.A(KEYINPUT43), .B(new_n906), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n851), .B1(new_n901), .B2(new_n904), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n906), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT44), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n921), .B(new_n906), .C1(new_n916), .C2(new_n917), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n893), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n918), .B2(new_n922), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT109), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n930), .A2(new_n933), .ZN(G397));
  NOR2_X1   g509(.A1(new_n491), .A2(new_n494), .ZN(new_n935));
  INV_X1    g510(.A(new_n487), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n468), .A2(new_n463), .ZN(new_n937));
  INV_X1    g512(.A(G138), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n471), .A2(new_n474), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(G1996), .A3(new_n745), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT112), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n732), .B(new_n738), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G1996), .B2(new_n745), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n794), .B(new_n789), .Z(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT111), .Z(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n947), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n935), .B2(new_n939), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n946), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G1971), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT113), .B1(G164), .B2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT50), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n946), .B1(new_n961), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(G2090), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(G8), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n976));
  INV_X1    g551(.A(G8), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(G166), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n979));
  NAND3_X1  g554(.A1(G303), .A2(G8), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n981), .ZN(new_n984));
  NAND2_X1  g559(.A1(G160), .A2(G40), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n972), .B2(new_n961), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n968), .A2(new_n970), .A3(KEYINPUT50), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n988), .A2(G2090), .B1(new_n966), .B2(G1971), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n989), .B2(G8), .ZN(new_n990));
  OR2_X1    g565(.A1(G305), .A2(G1981), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n586), .B1(new_n587), .B2(new_n509), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G1981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n968), .A2(new_n970), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n946), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n977), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n991), .A2(KEYINPUT49), .A3(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G288), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G1976), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n998), .A2(G8), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n983), .A2(new_n990), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1956), .B1(new_n986), .B2(new_n987), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n963), .A2(new_n965), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n574), .A2(new_n1017), .A3(new_n575), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(G299), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(new_n618), .A3(new_n1021), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  OR4_X1    g603(.A1(KEYINPUT122), .A2(new_n1013), .A3(new_n1016), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n988), .A2(new_n754), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n966), .A2(new_n1014), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT61), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(KEYINPUT122), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(KEYINPUT119), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1024), .A2(new_n1027), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1036), .A2(new_n1040), .A3(KEYINPUT120), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT120), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1029), .B(new_n1035), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n998), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n985), .B1(KEYINPUT45), .B2(new_n961), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n1047));
  INV_X1    g622(.A(G1996), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n964), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n964), .A2(new_n962), .A3(new_n1048), .A4(new_n946), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT121), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1045), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n558), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT59), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1055), .A3(new_n558), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1028), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1033), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1054), .A2(new_n1056), .B1(new_n1058), .B2(new_n1034), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n999), .A2(new_n738), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n706), .B1(new_n971), .B2(new_n973), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n610), .A2(KEYINPUT123), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n610), .A2(KEYINPUT123), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .A4(KEYINPUT60), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1043), .A2(new_n1059), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n607), .A3(new_n855), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1033), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n964), .A2(new_n962), .A3(new_n726), .A4(new_n946), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1076), .A2(KEYINPUT124), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT124), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n693), .B1(new_n971), .B2(new_n973), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1046), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n726), .A2(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(G301), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n963), .B1(new_n943), .B2(new_n944), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(KEYINPUT53), .A3(new_n726), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT54), .B(new_n1085), .C1(new_n1089), .C2(G301), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1089), .B2(G171), .ZN(new_n1092));
  OAI21_X1  g667(.A(G171), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT125), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(G171), .C1(new_n1080), .C2(new_n1084), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1966), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT116), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n971), .A2(G2084), .A3(new_n973), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1082), .A2(new_n1103), .A3(new_n1099), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(G168), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT51), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(G286), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1075), .A2(new_n1098), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1106), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1105), .B2(G8), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1107), .B(new_n1116), .C1(new_n1106), .C2(new_n1110), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1097), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1012), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1010), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1002), .A2(new_n1007), .A3(KEYINPUT115), .A4(new_n1009), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1002), .A2(new_n1005), .A3(new_n1003), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n991), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(new_n983), .B1(new_n1000), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1109), .A2(G8), .A3(G168), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n975), .A2(new_n981), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n982), .A2(KEYINPUT63), .A3(new_n1128), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n1127), .A2(new_n1129), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT63), .B1(new_n1011), .B2(new_n1127), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n960), .B1(new_n1119), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n957), .A2(new_n947), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT48), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n955), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n794), .A2(new_n789), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n953), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n732), .A2(G2067), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n947), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n948), .A2(new_n1048), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT46), .ZN(new_n1142));
  INV_X1    g717(.A(new_n951), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n948), .B1(new_n745), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NOR3_X1   g721(.A1(new_n1136), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1133), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1133), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g727(.A1(G401), .A2(G229), .ZN(new_n1154));
  AND2_X1   g728(.A1(new_n847), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g729(.A1(G227), .A2(new_n461), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n1158));
  XNOR2_X1  g732(.A(new_n1157), .B(new_n1158), .ZN(G308));
  XNOR2_X1  g733(.A(new_n1157), .B(KEYINPUT127), .ZN(G225));
endmodule


