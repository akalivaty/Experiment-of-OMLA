

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U551 ( .A(n522), .B(n521), .ZN(n531) );
  AND2_X1 U552 ( .A1(n710), .A2(n709), .ZN(n517) );
  NAND2_X1 U553 ( .A1(n700), .A2(n931), .ZN(n518) );
  AND2_X1 U554 ( .A1(n928), .A2(n755), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n742), .A2(n519), .ZN(n520) );
  AND2_X1 U556 ( .A1(n675), .A2(n673), .ZN(n662) );
  NOR2_X2 U557 ( .A1(n597), .A2(n711), .ZN(n648) );
  INV_X1 U558 ( .A(KEYINPUT106), .ZN(n698) );
  XNOR2_X1 U559 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U560 ( .A1(G543), .A2(n545), .ZN(n539) );
  AND2_X1 U561 ( .A1(n526), .A2(G2104), .ZN(n868) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n793) );
  NOR2_X1 U563 ( .A1(n579), .A2(G651), .ZN(n783) );
  NOR2_X1 U564 ( .A1(n630), .A2(n629), .ZN(n924) );
  NOR2_X1 U565 ( .A1(n538), .A2(n537), .ZN(G160) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U567 ( .A1(n871), .A2(G114), .ZN(n525) );
  XNOR2_X1 U568 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n531), .A2(G138), .ZN(n523) );
  XOR2_X1 U571 ( .A(KEYINPUT87), .B(n523), .Z(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n530) );
  INV_X1 U573 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U574 ( .A1(G102), .A2(n868), .ZN(n528) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n526), .ZN(n873) );
  NAND2_X1 U576 ( .A1(G126), .A2(n873), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U578 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U579 ( .A1(n531), .A2(G137), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G101), .A2(n868), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n532), .Z(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U583 ( .A1(G113), .A2(n871), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G125), .A2(n873), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U586 ( .A(G651), .ZN(n545) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n539), .Z(n785) );
  NAND2_X1 U588 ( .A1(G65), .A2(n785), .ZN(n541) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n579) );
  NAND2_X1 U590 ( .A1(G53), .A2(n783), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n793), .A2(G91), .ZN(n542) );
  XOR2_X1 U593 ( .A(KEYINPUT68), .B(n542), .Z(n543) );
  NOR2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X1 U595 ( .A1(n579), .A2(n545), .ZN(n789) );
  NAND2_X1 U596 ( .A1(n789), .A2(G78), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(G299) );
  NAND2_X1 U598 ( .A1(G64), .A2(n785), .ZN(n548) );
  XNOR2_X1 U599 ( .A(n548), .B(KEYINPUT67), .ZN(n553) );
  NAND2_X1 U600 ( .A1(G90), .A2(n793), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G77), .A2(n789), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U604 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n783), .A2(G52), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(G301) );
  INV_X1 U607 ( .A(G301), .ZN(G171) );
  NAND2_X1 U608 ( .A1(G63), .A2(n785), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G51), .A2(n783), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U611 ( .A(KEYINPUT6), .B(n558), .ZN(n565) );
  NAND2_X1 U612 ( .A1(n793), .A2(G89), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G76), .A2(n789), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT5), .B(n562), .ZN(n563) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(n563), .ZN(n564) );
  NOR2_X1 U618 ( .A1(n565), .A2(n564), .ZN(n567) );
  XOR2_X1 U619 ( .A(KEYINPUT74), .B(KEYINPUT7), .Z(n566) );
  XNOR2_X1 U620 ( .A(n567), .B(n566), .ZN(G168) );
  NAND2_X1 U621 ( .A1(G88), .A2(n793), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G75), .A2(n789), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U624 ( .A1(G62), .A2(n785), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G50), .A2(n783), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U627 ( .A1(n573), .A2(n572), .ZN(G166) );
  INV_X1 U628 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U629 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n574) );
  XNOR2_X1 U630 ( .A(n574), .B(G168), .ZN(G286) );
  NAND2_X1 U631 ( .A1(G49), .A2(n783), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n785), .A2(n577), .ZN(n578) );
  XOR2_X1 U635 ( .A(KEYINPUT83), .B(n578), .Z(n581) );
  NAND2_X1 U636 ( .A1(n579), .A2(G87), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(G288) );
  XOR2_X1 U638 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n583) );
  NAND2_X1 U639 ( .A1(G73), .A2(n789), .ZN(n582) );
  XNOR2_X1 U640 ( .A(n583), .B(n582), .ZN(n587) );
  NAND2_X1 U641 ( .A1(G61), .A2(n785), .ZN(n585) );
  NAND2_X1 U642 ( .A1(G48), .A2(n783), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U644 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n793), .A2(G86), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n589), .A2(n588), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G85), .A2(n793), .ZN(n591) );
  NAND2_X1 U648 ( .A1(G72), .A2(n789), .ZN(n590) );
  NAND2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U650 ( .A(KEYINPUT66), .B(n592), .Z(n596) );
  NAND2_X1 U651 ( .A1(G60), .A2(n785), .ZN(n594) );
  NAND2_X1 U652 ( .A1(G47), .A2(n783), .ZN(n593) );
  AND2_X1 U653 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U655 ( .A1(G164), .A2(G1384), .ZN(n712) );
  INV_X1 U656 ( .A(n712), .ZN(n597) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n711) );
  INV_X1 U658 ( .A(n648), .ZN(n667) );
  NAND2_X1 U659 ( .A1(n667), .A2(G8), .ZN(n708) );
  NOR2_X1 U660 ( .A1(G1966), .A2(n708), .ZN(n663) );
  XOR2_X1 U661 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n602) );
  NAND2_X1 U662 ( .A1(n648), .A2(G2072), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT27), .B(n598), .Z(n600) );
  NAND2_X1 U664 ( .A1(G1956), .A2(n667), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n638) );
  NAND2_X1 U666 ( .A1(n638), .A2(G299), .ZN(n601) );
  XOR2_X1 U667 ( .A(n602), .B(n601), .Z(n643) );
  XOR2_X1 U668 ( .A(G1996), .B(KEYINPUT97), .Z(n976) );
  NAND2_X1 U669 ( .A1(n976), .A2(n648), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT26), .ZN(n604) );
  XNOR2_X1 U671 ( .A(n604), .B(KEYINPUT64), .ZN(n618) );
  NAND2_X1 U672 ( .A1(n667), .A2(G1348), .ZN(n606) );
  INV_X1 U673 ( .A(KEYINPUT99), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G2067), .A2(n648), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n634) );
  NAND2_X1 U677 ( .A1(G92), .A2(n793), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G66), .A2(n785), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U680 ( .A1(G79), .A2(n789), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G54), .A2(n783), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(KEYINPUT72), .B(n613), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n616), .B(KEYINPUT15), .ZN(n915) );
  NAND2_X1 U686 ( .A1(n634), .A2(n915), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n633) );
  NAND2_X1 U688 ( .A1(n667), .A2(G1341), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT98), .ZN(n631) );
  NAND2_X1 U690 ( .A1(G56), .A2(n785), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT70), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT14), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G43), .A2(n783), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n630) );
  NAND2_X1 U695 ( .A1(n793), .A2(G81), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(KEYINPUT12), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G68), .A2(n789), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U699 ( .A(KEYINPUT13), .B(n627), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT71), .B(n628), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n631), .A2(n924), .ZN(n632) );
  NOR2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n636) );
  NOR2_X1 U703 ( .A1(n634), .A2(n915), .ZN(n635) );
  NOR2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U705 ( .A(KEYINPUT100), .B(n637), .ZN(n640) );
  OR2_X1 U706 ( .A1(G299), .A2(n638), .ZN(n639) );
  AND2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U708 ( .A(n641), .B(KEYINPUT101), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n643), .A2(n642), .ZN(n645) );
  INV_X1 U710 ( .A(KEYINPUT29), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n653) );
  NOR2_X1 U712 ( .A1(n648), .A2(G1961), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(KEYINPUT93), .ZN(n650) );
  XNOR2_X1 U714 ( .A(G2078), .B(KEYINPUT25), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT94), .ZN(n970) );
  NAND2_X1 U716 ( .A1(n970), .A2(n648), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n655) );
  AND2_X1 U718 ( .A1(n655), .A2(G171), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT95), .B(n651), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U721 ( .A(KEYINPUT102), .B(n654), .ZN(n675) );
  NOR2_X1 U722 ( .A1(G171), .A2(n655), .ZN(n660) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n667), .ZN(n664) );
  NOR2_X1 U724 ( .A1(n663), .A2(n664), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G8), .A2(n656), .ZN(n657) );
  XNOR2_X1 U726 ( .A(KEYINPUT30), .B(n657), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n658), .A2(G168), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U729 ( .A(KEYINPUT31), .B(n661), .Z(n673) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U731 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n683) );
  INV_X1 U733 ( .A(G8), .ZN(n672) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n708), .ZN(n669) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n670), .A2(G303), .ZN(n671) );
  OR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n676) );
  AND2_X1 U739 ( .A1(n673), .A2(n676), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n679) );
  INV_X1 U741 ( .A(n676), .ZN(n677) );
  OR2_X1 U742 ( .A1(n677), .A2(G286), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n681) );
  XOR2_X1 U744 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n703) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U748 ( .A1(G288), .A2(G1976), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT104), .ZN(n913) );
  NOR2_X1 U750 ( .A1(n685), .A2(n913), .ZN(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT105), .B(n686), .Z(n688) );
  INV_X1 U752 ( .A(n708), .ZN(n692) );
  NAND2_X1 U753 ( .A1(n913), .A2(n692), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n687), .A2(KEYINPUT33), .ZN(n690) );
  AND2_X1 U755 ( .A1(n688), .A2(n690), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n703), .A2(n689), .ZN(n697) );
  INV_X1 U757 ( .A(n690), .ZN(n695) );
  INV_X1 U758 ( .A(KEYINPUT33), .ZN(n691) );
  NAND2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n925) );
  AND2_X1 U760 ( .A1(n691), .A2(n925), .ZN(n693) );
  AND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n699) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n931) );
  NAND2_X1 U765 ( .A1(G8), .A2(G166), .ZN(n701) );
  NOR2_X1 U766 ( .A1(G2090), .A2(n701), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(KEYINPUT107), .ZN(n704) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U769 ( .A1(n705), .A2(n708), .ZN(n710) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U771 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  OR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n518), .A2(n517), .ZN(n743) );
  NOR2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n755) );
  NAND2_X1 U775 ( .A1(G140), .A2(n531), .ZN(n714) );
  NAND2_X1 U776 ( .A1(G104), .A2(n868), .ZN(n713) );
  NAND2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U778 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U779 ( .A1(G116), .A2(n871), .ZN(n717) );
  NAND2_X1 U780 ( .A1(G128), .A2(n873), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U782 ( .A(n718), .B(KEYINPUT35), .Z(n719) );
  NOR2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U784 ( .A(KEYINPUT36), .B(n721), .Z(n722) );
  XOR2_X1 U785 ( .A(KEYINPUT88), .B(n722), .Z(n879) );
  XNOR2_X1 U786 ( .A(KEYINPUT37), .B(G2067), .ZN(n752) );
  NOR2_X1 U787 ( .A1(n879), .A2(n752), .ZN(n1009) );
  NAND2_X1 U788 ( .A1(n755), .A2(n1009), .ZN(n750) );
  NAND2_X1 U789 ( .A1(n873), .A2(G129), .ZN(n729) );
  NAND2_X1 U790 ( .A1(G141), .A2(n531), .ZN(n724) );
  NAND2_X1 U791 ( .A1(G117), .A2(n871), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n868), .A2(G105), .ZN(n725) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n725), .Z(n726) );
  NOR2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U797 ( .A(KEYINPUT91), .B(n730), .Z(n887) );
  NAND2_X1 U798 ( .A1(n887), .A2(G1996), .ZN(n740) );
  NAND2_X1 U799 ( .A1(G95), .A2(n868), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n731), .B(KEYINPUT90), .ZN(n738) );
  NAND2_X1 U801 ( .A1(G131), .A2(n531), .ZN(n733) );
  NAND2_X1 U802 ( .A1(G119), .A2(n873), .ZN(n732) );
  NAND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U804 ( .A1(G107), .A2(n871), .ZN(n734) );
  XNOR2_X1 U805 ( .A(KEYINPUT89), .B(n734), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n856) );
  NAND2_X1 U808 ( .A1(n856), .A2(G1991), .ZN(n739) );
  NAND2_X1 U809 ( .A1(n740), .A2(n739), .ZN(n992) );
  NAND2_X1 U810 ( .A1(n992), .A2(n755), .ZN(n744) );
  NAND2_X1 U811 ( .A1(n750), .A2(n744), .ZN(n741) );
  XNOR2_X1 U812 ( .A(n741), .B(KEYINPUT92), .ZN(n742) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n928) );
  NAND2_X1 U814 ( .A1(n743), .A2(n520), .ZN(n758) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n887), .ZN(n1006) );
  INV_X1 U816 ( .A(n744), .ZN(n747) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n856), .ZN(n996) );
  NOR2_X1 U819 ( .A1(n745), .A2(n996), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n1006), .A2(n748), .ZN(n749) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n749), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n879), .A2(n752), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT108), .ZN(n1015) );
  NAND2_X1 U826 ( .A1(n754), .A2(n1015), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U829 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U831 ( .A(G57), .ZN(G237) );
  INV_X1 U832 ( .A(G132), .ZN(G219) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U835 ( .A(n760), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U836 ( .A(G223), .B(KEYINPUT69), .ZN(n825) );
  NAND2_X1 U837 ( .A1(n825), .A2(G567), .ZN(n761) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  NAND2_X1 U839 ( .A1(n924), .A2(G860), .ZN(G153) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n763) );
  INV_X1 U841 ( .A(G868), .ZN(n799) );
  NAND2_X1 U842 ( .A1(n915), .A2(n799), .ZN(n762) );
  NAND2_X1 U843 ( .A1(n763), .A2(n762), .ZN(G284) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n764) );
  XNOR2_X1 U845 ( .A(n764), .B(KEYINPUT76), .ZN(n766) );
  NOR2_X1 U846 ( .A1(G286), .A2(n799), .ZN(n765) );
  NOR2_X1 U847 ( .A1(n766), .A2(n765), .ZN(G297) );
  INV_X1 U848 ( .A(G860), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n767), .A2(G559), .ZN(n768) );
  INV_X1 U850 ( .A(n915), .ZN(n892) );
  NAND2_X1 U851 ( .A1(n768), .A2(n892), .ZN(n769) );
  XNOR2_X1 U852 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U853 ( .A1(n892), .A2(G868), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G559), .A2(n770), .ZN(n772) );
  AND2_X1 U855 ( .A1(n799), .A2(n924), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(G282) );
  XOR2_X1 U857 ( .A(G2100), .B(KEYINPUT78), .Z(n782) );
  NAND2_X1 U858 ( .A1(G135), .A2(n531), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G111), .A2(n871), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n873), .A2(G123), .ZN(n775) );
  XOR2_X1 U862 ( .A(KEYINPUT18), .B(n775), .Z(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n868), .A2(G99), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n993) );
  XNOR2_X1 U866 ( .A(KEYINPUT77), .B(n993), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(G2096), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U869 ( .A1(n783), .A2(G55), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT81), .B(n784), .Z(n787) );
  NAND2_X1 U871 ( .A1(n785), .A2(G67), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U873 ( .A(KEYINPUT82), .B(n788), .ZN(n792) );
  NAND2_X1 U874 ( .A1(n789), .A2(G80), .ZN(n790) );
  XOR2_X1 U875 ( .A(KEYINPUT80), .B(n790), .Z(n791) );
  NOR2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U877 ( .A1(n793), .A2(G93), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n808) );
  NAND2_X1 U879 ( .A1(G559), .A2(n892), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT79), .ZN(n809) );
  XNOR2_X1 U881 ( .A(n924), .B(n809), .ZN(n797) );
  NOR2_X1 U882 ( .A1(G860), .A2(n797), .ZN(n798) );
  XOR2_X1 U883 ( .A(n808), .B(n798), .Z(G145) );
  NAND2_X1 U884 ( .A1(n799), .A2(n808), .ZN(n800) );
  XNOR2_X1 U885 ( .A(n800), .B(KEYINPUT86), .ZN(n812) );
  XNOR2_X1 U886 ( .A(KEYINPUT19), .B(G299), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(G288), .ZN(n802) );
  XNOR2_X1 U888 ( .A(KEYINPUT85), .B(n802), .ZN(n804) );
  XNOR2_X1 U889 ( .A(G290), .B(n924), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n804), .B(n803), .ZN(n805) );
  XNOR2_X1 U891 ( .A(G166), .B(n805), .ZN(n806) );
  XNOR2_X1 U892 ( .A(n806), .B(G305), .ZN(n807) );
  XOR2_X1 U893 ( .A(n808), .B(n807), .Z(n891) );
  XNOR2_X1 U894 ( .A(n891), .B(n809), .ZN(n810) );
  NAND2_X1 U895 ( .A1(G868), .A2(n810), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n817) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n817), .Z(n818) );
  NOR2_X1 U905 ( .A1(G218), .A2(n818), .ZN(n819) );
  NAND2_X1 U906 ( .A1(G96), .A2(n819), .ZN(n829) );
  NAND2_X1 U907 ( .A1(n829), .A2(G2106), .ZN(n823) );
  NAND2_X1 U908 ( .A1(G120), .A2(G108), .ZN(n820) );
  NOR2_X1 U909 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U910 ( .A1(G69), .A2(n821), .ZN(n830) );
  NAND2_X1 U911 ( .A1(n830), .A2(G567), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n831) );
  NAND2_X1 U913 ( .A1(G483), .A2(G661), .ZN(n824) );
  NOR2_X1 U914 ( .A1(n831), .A2(n824), .ZN(n828) );
  NAND2_X1 U915 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n831), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2096), .B(G2100), .Z(n833) );
  XNOR2_X1 U929 ( .A(KEYINPUT42), .B(G2678), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2090), .Z(n835) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1966), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1956), .B(G1981), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1961), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U947 ( .A1(G124), .A2(n873), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n871), .A2(G112), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U951 ( .A1(G136), .A2(n531), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G100), .A2(n868), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(G162) );
  XNOR2_X1 U955 ( .A(G164), .B(n856), .ZN(n867) );
  NAND2_X1 U956 ( .A1(G142), .A2(n531), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G106), .A2(n868), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT45), .B(n859), .ZN(n865) );
  NAND2_X1 U960 ( .A1(G118), .A2(n871), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT111), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G130), .A2(n873), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT110), .B(n861), .Z(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n883) );
  NAND2_X1 U967 ( .A1(G139), .A2(n531), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G103), .A2(n868), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n878) );
  NAND2_X1 U970 ( .A1(n871), .A2(G115), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT112), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G127), .A2(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n1001) );
  XOR2_X1 U976 ( .A(G162), .B(n1001), .Z(n881) );
  XNOR2_X1 U977 ( .A(G160), .B(n879), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n889) );
  XNOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n993), .B(KEYINPUT113), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U985 ( .A1(G37), .A2(n890), .ZN(G395) );
  XOR2_X1 U986 ( .A(KEYINPUT114), .B(n891), .Z(n894) );
  XNOR2_X1 U987 ( .A(G171), .B(n892), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(n895), .B(G286), .Z(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2430), .B(G2451), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2446), .B(G2427), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n905) );
  XOR2_X1 U994 ( .A(G2438), .B(KEYINPUT109), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2443), .B(G2454), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n901), .B(G2435), .Z(n903) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(n906), .A2(G14), .ZN(n912) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(n912), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(G16), .B(KEYINPUT56), .ZN(n939) );
  XOR2_X1 U1012 ( .A(n913), .B(KEYINPUT125), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1961), .B(KEYINPUT122), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(G301), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(G1348), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(KEYINPUT123), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n937) );
  XNOR2_X1 U1019 ( .A(G1956), .B(KEYINPUT124), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n921), .B(G299), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G1971), .B(G303), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(n924), .B(G1341), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT57), .B(n933), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n965) );
  INV_X1 U1033 ( .A(G16), .ZN(n963) );
  XOR2_X1 U1034 ( .A(G1348), .B(KEYINPUT59), .Z(n940) );
  XNOR2_X1 U1035 ( .A(G4), .B(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(G20), .B(G1956), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G6), .B(G1981), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT126), .B(n947), .Z(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT60), .B(n948), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G21), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G5), .B(G1961), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G24), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G1971), .B(KEYINPUT127), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(n955), .B(G22), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT58), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT61), .B(n961), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G2084), .B(G34), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT54), .ZN(n984) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1062 ( .A(G1991), .B(G25), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G2067), .B(G26), .Z(n969) );
  NAND2_X1 U1066 ( .A1(n969), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G27), .B(n970), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT119), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G32), .B(n976), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT120), .B(n982), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT55), .B(n985), .ZN(n987) );
  INV_X1 U1078 ( .A(G29), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n988), .A2(G11), .ZN(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT121), .B(n989), .Z(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n1022) );
  INV_X1 U1083 ( .A(KEYINPUT55), .ZN(n1018) );
  INV_X1 U1084 ( .A(n992), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G160), .B(G2084), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT116), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1013) );
  XNOR2_X1 U1090 ( .A(G164), .B(G2078), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT117), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1001), .Z(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1004), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT51), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .Z(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1020), .B(KEYINPUT118), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

