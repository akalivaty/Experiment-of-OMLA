//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT65), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT65), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AOI211_X1 g019(.A(KEYINPUT64), .B(new_n199), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(G143), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(new_n210), .B2(G143), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n201), .A3(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n206), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n199), .B1(new_n203), .B2(new_n205), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n219), .B2(KEYINPUT64), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n198), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n188), .A2(G137), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT67), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n190), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(G131), .C1(new_n225), .C2(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n196), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT65), .B(G146), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G143), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n207), .A2(new_n208), .A3(G143), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n230), .A2(new_n231), .B1(new_n204), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n209), .A2(new_n211), .A3(new_n213), .A4(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n227), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n238), .A2(KEYINPUT30), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(KEYINPUT30), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n221), .A2(new_n237), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(new_n199), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n242), .B(new_n243), .C1(new_n232), .C2(new_n204), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n216), .A3(new_n214), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT64), .B(new_n243), .C1(new_n232), .C2(new_n204), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n215), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n197), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n238), .B(KEYINPUT30), .C1(new_n248), .C2(new_n236), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G116), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G119), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n255), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n259), .A2(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n248), .A2(new_n261), .A3(new_n236), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT26), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G101), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT26), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n269), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G101), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n262), .A2(new_n264), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n275), .A3(KEYINPUT70), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n261), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n221), .B2(new_n237), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n285), .B2(new_n263), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n263), .A2(KEYINPUT28), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n263), .B1(new_n250), .B2(new_n261), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n277), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n279), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G472), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n290), .A2(new_n277), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n287), .A2(new_n286), .ZN(new_n301));
  INV_X1    g115(.A(new_n283), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n287), .A2(new_n286), .A3(KEYINPUT29), .A4(new_n277), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G472), .B1(new_n305), .B2(G902), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n294), .A4(new_n295), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n298), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G952), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(G234), .A2(G237), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT21), .B(G898), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(G902), .A3(G953), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT86), .B1(new_n201), .B2(G128), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT86), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n231), .A3(G143), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n201), .A2(G128), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n323), .A2(KEYINPUT88), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT88), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(new_n188), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n231), .B2(G143), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n201), .A2(KEYINPUT86), .A3(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(KEYINPUT88), .A3(new_n324), .ZN(new_n333));
  AOI21_X1  g147(.A(G134), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT89), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G107), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT85), .A2(G122), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT85), .A2(G122), .ZN(new_n338));
  OAI21_X1  g152(.A(G116), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n336), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g154(.A(G122), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(G116), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n188), .B1(new_n325), .B2(new_n326), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(G134), .A3(new_n333), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n340), .A2(new_n342), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n335), .A2(new_n343), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n324), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT87), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n323), .B1(KEYINPUT13), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g167(.A(G134), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n342), .B(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n344), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(KEYINPUT9), .B(G234), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G217), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(G953), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n349), .A2(new_n356), .A3(new_n361), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT90), .ZN(new_n366));
  INV_X1    g180(.A(G478), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT15), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n349), .A2(new_n356), .A3(new_n361), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n361), .B1(new_n349), .B2(new_n356), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n366), .B(new_n295), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n368), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  INV_X1    g190(.A(G125), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n229), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT16), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n375), .A3(G125), .ZN(new_n384));
  OAI211_X1 g198(.A(G146), .B(new_n384), .C1(new_n379), .C2(new_n383), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n201), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n201), .A2(KEYINPUT84), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(G214), .A3(new_n265), .A4(new_n266), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n195), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n195), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n382), .B(new_n385), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n376), .A2(new_n378), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n229), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n210), .B2(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n387), .B(new_n389), .C1(new_n397), .C2(new_n195), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n387), .A2(new_n389), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G131), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n396), .B(new_n398), .C1(new_n400), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT17), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n408), .A3(new_n391), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n384), .B1(new_n379), .B2(new_n383), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n210), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(KEYINPUT17), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n409), .A2(new_n385), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n405), .A3(new_n401), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G475), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n295), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n420), .A3(new_n416), .A4(new_n295), .ZN(new_n421));
  INV_X1    g235(.A(new_n414), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n405), .B1(new_n413), .B2(new_n401), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n295), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n419), .A2(new_n421), .B1(G475), .B2(new_n424), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n319), .A2(new_n370), .A3(new_n374), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G469), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT3), .B1(new_n404), .B2(G107), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT3), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n336), .A3(G104), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n404), .A2(G107), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n274), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n336), .A2(G104), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n404), .A2(G107), .ZN(new_n435));
  OAI21_X1  g249(.A(G101), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G128), .B1(new_n204), .B2(new_n228), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n214), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n439), .B2(new_n235), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT76), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n442), .B(new_n437), .C1(new_n439), .C2(new_n235), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n428), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G101), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT4), .A3(new_n433), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n448), .A3(G101), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n245), .A2(new_n247), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n437), .B1(new_n233), .B2(new_n235), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n451), .A2(new_n452), .B1(new_n453), .B2(KEYINPUT10), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n444), .A2(new_n197), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(G110), .B(G140), .Z(new_n456));
  AND2_X1   g270(.A1(new_n266), .A2(G227), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n233), .A2(new_n235), .ZN(new_n460));
  INV_X1    g274(.A(new_n437), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n441), .A2(new_n443), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT77), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n462), .B(new_n198), .C1(new_n463), .C2(KEYINPUT12), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n198), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n198), .B2(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n459), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n444), .A2(new_n454), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n198), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n458), .B1(new_n470), .B2(new_n455), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n427), .B(new_n295), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n455), .A3(new_n458), .ZN(new_n473));
  INV_X1    g287(.A(new_n455), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n464), .B2(new_n467), .ZN(new_n475));
  OAI211_X1 g289(.A(G469), .B(new_n473), .C1(new_n475), .C2(new_n458), .ZN(new_n476));
  NAND2_X1  g290(.A1(G469), .A2(G902), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n359), .B2(G902), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n426), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n360), .B1(G234), .B2(new_n295), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n231), .A2(G119), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT23), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n252), .B2(G128), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n484), .B(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT71), .B1(new_n252), .B2(G128), .ZN(new_n488));
  MUX2_X1   g302(.A(KEYINPUT71), .B(new_n488), .S(new_n483), .Z(new_n489));
  XOR2_X1   g303(.A(KEYINPUT24), .B(G110), .Z(new_n490));
  OAI22_X1  g304(.A1(new_n487), .A2(G110), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n385), .A3(new_n395), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n411), .A2(new_n385), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(G110), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n490), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n491), .A2(new_n498), .A3(new_n385), .A4(new_n395), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT22), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(G137), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n493), .A2(new_n497), .A3(new_n499), .A4(new_n503), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n295), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n505), .A2(KEYINPUT25), .A3(new_n295), .A4(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n482), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n505), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n505), .B2(new_n506), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n481), .A2(G902), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT75), .Z(new_n516));
  NOR3_X1   g330(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n245), .A2(G125), .A3(new_n247), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n231), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n207), .A2(new_n208), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n204), .B1(new_n524), .B2(new_n201), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n377), .B(new_n235), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n521), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n521), .ZN(new_n529));
  INV_X1    g343(.A(G224), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n528), .A2(KEYINPUT7), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT81), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n534), .B2(KEYINPUT7), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n534), .B2(KEYINPUT7), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n210), .A2(KEYINPUT66), .A3(G143), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n229), .B2(G143), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n215), .B1(new_n538), .B2(new_n211), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n539), .A2(new_n244), .B1(new_n246), .B2(new_n215), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT79), .B1(new_n540), .B2(G125), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n527), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G113), .B1(new_n253), .B2(KEYINPUT5), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT5), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n259), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n260), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n461), .ZN(new_n547));
  XOR2_X1   g361(.A(G110), .B(G122), .Z(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT8), .Z(new_n549));
  NOR3_X1   g363(.A1(new_n256), .A2(new_n257), .A3(new_n544), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n260), .B1(new_n550), .B2(new_n543), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n547), .B(new_n549), .C1(new_n551), .C2(new_n461), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n261), .A2(new_n449), .A3(new_n447), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n461), .B(new_n260), .C1(new_n550), .C2(new_n543), .ZN(new_n554));
  INV_X1    g368(.A(new_n548), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n533), .A2(new_n542), .A3(new_n552), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n531), .B1(new_n527), .B2(new_n541), .ZN(new_n558));
  INV_X1    g372(.A(new_n526), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n540), .B2(G125), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n529), .B(new_n532), .C1(new_n560), .C2(new_n521), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT80), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT80), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n553), .A2(new_n555), .A3(new_n554), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n555), .B1(new_n553), .B2(new_n554), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n553), .A2(new_n554), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n548), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT6), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT78), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n556), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n295), .B(new_n557), .C1(new_n564), .C2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G210), .B1(G237), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n572), .B(new_n575), .C1(new_n562), .C2(new_n563), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(new_n295), .A3(new_n580), .A4(new_n557), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n520), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n308), .A2(new_n480), .A3(new_n518), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AOI21_X1  g401(.A(new_n291), .B1(new_n290), .B2(new_n277), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n284), .B1(new_n241), .B2(new_n249), .ZN(new_n589));
  NOR4_X1   g403(.A1(new_n589), .A2(KEYINPUT31), .A3(new_n263), .A4(new_n276), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n588), .A2(new_n590), .A3(new_n288), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n591), .B2(G902), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n592), .A2(new_n296), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n478), .A2(new_n518), .A3(new_n479), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n577), .A2(new_n578), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n583), .A2(new_n295), .A3(new_n579), .A4(new_n557), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n519), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n597), .A2(KEYINPUT92), .A3(new_n519), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n318), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n371), .A2(new_n372), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT33), .B1(new_n372), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n363), .B(new_n364), .C1(KEYINPUT93), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(G478), .B(new_n295), .C1(new_n608), .C2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n365), .A2(G478), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n425), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n604), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n596), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND2_X1  g433(.A1(new_n370), .A2(new_n374), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n424), .A2(G475), .ZN(new_n622));
  INV_X1    g436(.A(new_n419), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n417), .A2(new_n418), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n604), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n596), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(new_n511), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n504), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n500), .B(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n516), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n480), .A2(new_n593), .A3(new_n585), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT37), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G110), .ZN(G12));
  NAND2_X1  g453(.A1(new_n308), .A2(new_n636), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n601), .A2(new_n602), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n478), .A2(new_n479), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n317), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n312), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n622), .B(new_n646), .C1(new_n623), .C2(new_n624), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n621), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  AND2_X1   g464(.A1(new_n582), .A2(new_n584), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT38), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n652), .A2(new_n520), .A3(new_n621), .A4(new_n425), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n302), .B1(new_n263), .B2(new_n285), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n278), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n655), .B2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n298), .A2(new_n307), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n478), .A2(new_n479), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n646), .B(KEYINPUT39), .Z(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n636), .B1(new_n661), .B2(KEYINPUT40), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n653), .A2(new_n657), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NAND2_X1  g479(.A1(new_n612), .A2(new_n614), .ZN(new_n666));
  INV_X1    g480(.A(new_n425), .ZN(new_n667));
  AND4_X1   g481(.A1(KEYINPUT94), .A2(new_n666), .A3(new_n667), .A4(new_n646), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT94), .B1(new_n615), .B2(new_n646), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n641), .A3(new_n642), .A4(new_n643), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NAND2_X1  g486(.A1(new_n308), .A2(new_n518), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n468), .A2(new_n471), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n427), .B1(new_n674), .B2(new_n295), .ZN(new_n675));
  INV_X1    g489(.A(new_n472), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n479), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n616), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT41), .B(G113), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NOR2_X1   g497(.A1(new_n627), .A2(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n254), .ZN(G18));
  AND2_X1   g499(.A1(new_n677), .A2(new_n479), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n641), .A2(new_n642), .A3(new_n426), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NAND3_X1  g502(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n296), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT95), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n293), .A2(new_n690), .A3(new_n294), .A4(new_n295), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n686), .A2(new_n692), .A3(new_n518), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n621), .A2(new_n425), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n604), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  AOI22_X1  g510(.A1(new_n689), .A2(new_n691), .B1(new_n631), .B2(new_n635), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n670), .A2(new_n642), .A3(new_n686), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  AND3_X1   g513(.A1(new_n582), .A2(new_n519), .A3(new_n584), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n643), .A3(KEYINPUT96), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT96), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n582), .A2(new_n519), .A3(new_n584), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n658), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n701), .A2(new_n704), .A3(new_n518), .A4(new_n308), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n670), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n363), .A2(new_n364), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n363), .A2(KEYINPUT93), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT33), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n367), .B(G902), .C1(new_n711), .C2(new_n610), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n667), .B(new_n646), .C1(new_n712), .C2(new_n613), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT94), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n615), .A2(KEYINPUT94), .A3(new_n646), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n708), .B1(new_n705), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n707), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n195), .ZN(G33));
  INV_X1    g535(.A(new_n673), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n648), .A3(new_n704), .A4(new_n701), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  AOI21_X1  g538(.A(new_n667), .B1(new_n612), .B2(new_n614), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT43), .ZN(new_n726));
  INV_X1    g540(.A(new_n593), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n636), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n700), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT98), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n473), .B1(new_n475), .B2(new_n458), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n739), .B2(new_n477), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n676), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n477), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n479), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n659), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n730), .A2(KEYINPUT98), .A3(new_n700), .A4(new_n731), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n734), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  AND2_X1   g562(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR4_X1    g565(.A1(new_n518), .A2(new_n717), .A3(new_n308), .A4(new_n703), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT99), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n726), .A2(new_n313), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n693), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n642), .ZN(new_n761));
  INV_X1    g575(.A(new_n615), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n657), .A2(new_n312), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n518), .A3(new_n686), .A4(new_n700), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n761), .B(new_n310), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n759), .A2(new_n700), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n680), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT113), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n770), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n775), .A3(new_n770), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n771), .A2(new_n772), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n758), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n760), .A2(new_n520), .A3(new_n652), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n760), .A2(KEYINPUT50), .A3(new_n520), .A4(new_n652), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n768), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n686), .A3(new_n697), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n764), .A2(new_n667), .A3(new_n666), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n677), .B(KEYINPUT101), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n749), .A2(new_n750), .B1(new_n479), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n518), .A3(new_n692), .A4(new_n784), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n787), .B(new_n791), .C1(new_n792), .C2(KEYINPUT51), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n783), .A3(new_n785), .A4(new_n786), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n783), .A2(new_n792), .A3(new_n785), .A4(new_n786), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n778), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n767), .A2(new_n777), .A3(new_n758), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n601), .A2(new_n643), .A3(new_n602), .A4(new_n694), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n646), .B(KEYINPUT107), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n636), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n657), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n671), .A2(new_n698), .A3(new_n649), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT108), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n800), .A2(new_n803), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n640), .A2(new_n603), .A3(new_n658), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n670), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n649), .A4(new_n698), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n648), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n715), .A2(new_n692), .A3(new_n636), .A4(new_n716), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n701), .A2(new_n704), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n705), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n703), .A2(new_n658), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n620), .A2(new_n647), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n641), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT105), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n815), .A2(new_n816), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT105), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n723), .A3(new_n824), .A4(new_n820), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(new_n719), .A3(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n679), .B(new_n604), .C1(new_n615), .C2(new_n626), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n695), .A3(new_n687), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n520), .B(new_n318), .C1(new_n582), .C2(new_n584), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n369), .B1(new_n365), .B2(new_n366), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n373), .A2(new_n368), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n425), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT102), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n620), .A2(KEYINPUT102), .A3(new_n425), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n829), .A2(new_n593), .A3(new_n594), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n637), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT103), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n829), .A2(new_n615), .A3(new_n593), .A4(new_n594), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n841), .A2(new_n586), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(new_n637), .A3(KEYINPUT103), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT104), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT104), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n846), .A3(new_n842), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n828), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n813), .A2(new_n826), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n698), .A2(new_n649), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT106), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n698), .A2(new_n649), .A3(KEYINPUT106), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n671), .A3(new_n804), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n698), .A2(new_n649), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n810), .B1(new_n858), .B2(new_n809), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n805), .A2(KEYINPUT108), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n813), .A3(new_n848), .A4(new_n826), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n812), .B1(new_n806), .B2(new_n811), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n849), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n862), .A2(KEYINPUT109), .A3(new_n863), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n798), .A2(new_n799), .A3(new_n865), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n309), .A2(new_n266), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n788), .B(KEYINPUT49), .ZN(new_n877));
  INV_X1    g691(.A(new_n657), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n725), .A2(new_n518), .A3(new_n519), .A4(new_n479), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT100), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n652), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT115), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(G75));
  AND3_X1   g700(.A1(new_n862), .A2(KEYINPUT109), .A3(new_n863), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT109), .B1(new_n862), .B2(new_n863), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n849), .A2(new_n855), .A3(new_n863), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n295), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n891), .B2(G210), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n564), .A2(new_n576), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n583), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  AOI211_X1 g711(.A(KEYINPUT56), .B(new_n895), .C1(new_n891), .C2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n266), .A2(G952), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G51));
  NAND3_X1  g714(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT54), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n901), .B2(KEYINPUT54), .ZN(new_n904));
  INV_X1    g718(.A(new_n873), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n477), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n674), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n739), .B(KEYINPUT118), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n891), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n909), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  INV_X1    g727(.A(new_n415), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n899), .ZN(G60));
  INV_X1    g731(.A(new_n899), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n873), .B2(new_n865), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n608), .A2(new_n611), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT119), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n906), .ZN(new_n925));
  INV_X1    g739(.A(new_n920), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(G63));
  NOR2_X1   g742(.A1(new_n513), .A2(new_n514), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n890), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(KEYINPUT121), .A3(new_n918), .ZN(new_n934));
  INV_X1    g748(.A(new_n932), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n901), .A2(new_n633), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n929), .B1(new_n901), .B2(new_n935), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n899), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n918), .A4(new_n936), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n315), .B2(new_n530), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n848), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n576), .B1(G898), .B2(new_n266), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  AND2_X1   g762(.A1(new_n852), .A2(new_n853), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n671), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n745), .A2(new_n722), .A3(new_n642), .A4(new_n694), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n951), .A2(new_n719), .A3(new_n723), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n952), .A3(new_n747), .A4(new_n756), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n266), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n644), .A2(G953), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n380), .A2(new_n381), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n250), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g776(.A(new_n960), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n949), .A2(new_n664), .A3(new_n671), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n747), .A2(new_n756), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n762), .A2(new_n834), .A3(new_n835), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n722), .A2(new_n660), .A3(new_n700), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n970), .B2(G953), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n958), .A2(new_n972), .A3(new_n960), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n962), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n971), .A2(new_n978), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n961), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n974), .A2(new_n983), .A3(new_n975), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n977), .A2(new_n982), .A3(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  NOR3_X1   g801(.A1(new_n589), .A2(new_n263), .A3(new_n276), .ZN(new_n988));
  OAI221_X1 g802(.A(new_n987), .B1(new_n299), .B2(new_n988), .C1(new_n857), .C2(new_n864), .ZN(new_n989));
  INV_X1    g803(.A(new_n848), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n953), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n290), .B(KEYINPUT127), .Z(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n276), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n918), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n970), .A2(new_n848), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n987), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT126), .B1(new_n995), .B2(new_n987), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n996), .A2(new_n997), .A3(new_n992), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n998), .B2(new_n277), .ZN(G57));
endmodule


