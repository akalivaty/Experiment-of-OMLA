//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT26), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  AND2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G183gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(new_n217), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT28), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n214), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(new_n213), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n218), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G176gat), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n207), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n212), .B2(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(G183gat), .B(G190gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n241), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n232), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n243), .A2(new_n241), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n232), .B1(new_n234), .B2(new_n206), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n246), .A2(new_n242), .A3(new_n239), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT68), .B(G120gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n254), .B(new_n257), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n256), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g060(.A1(G113gat), .A2(G120gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(new_n253), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n231), .A2(new_n249), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n259), .B(new_n271), .C1(new_n266), .C2(new_n267), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n231), .A2(new_n249), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n205), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G15gat), .B(G43gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n226), .A2(new_n230), .B1(new_n245), .B2(new_n248), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n269), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n269), .A2(new_n272), .ZN(new_n284));
  OAI221_X1 g083(.A(new_n283), .B1(new_n202), .B2(new_n203), .C1(new_n284), .C2(new_n282), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n270), .A2(new_n273), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n205), .A2(KEYINPUT34), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n285), .A2(KEYINPUT34), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n280), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n274), .B(KEYINPUT32), .C1(new_n276), .C2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n281), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n281), .B2(new_n290), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n281), .A2(new_n290), .ZN(new_n294));
  INV_X1    g093(.A(new_n288), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n288), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n298));
  OR2_X1    g097(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n308));
  OAI21_X1  g107(.A(G218gat), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310));
  AOI221_X4 g109(.A(KEYINPUT73), .B1(new_n305), .B2(new_n306), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n306), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n304), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT72), .B(G211gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT22), .B1(new_n317), .B2(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n314), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT73), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n312), .A3(new_n314), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n303), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n229), .B1(new_n228), .B2(new_n218), .ZN(new_n325));
  AND4_X1   g124(.A1(new_n216), .A2(new_n220), .A3(new_n222), .A4(new_n217), .ZN(new_n326));
  NOR4_X1   g125(.A1(new_n227), .A2(new_n326), .A3(new_n213), .A4(KEYINPUT66), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n249), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n231), .A2(KEYINPUT75), .A3(new_n249), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT74), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n249), .A2(new_n225), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n324), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n231), .A2(KEYINPUT75), .A3(new_n249), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT75), .B1(new_n231), .B2(new_n249), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(new_n331), .A3(new_n336), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n323), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR4_X1   g152(.A1(new_n342), .A2(new_n347), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n336), .B1(new_n330), .B2(new_n332), .ZN(new_n355));
  INV_X1    g154(.A(new_n346), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n324), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n340), .B1(new_n333), .B2(new_n336), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n357), .B(new_n350), .C1(new_n358), .C2(new_n324), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n357), .B1(new_n358), .B2(new_n324), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n351), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n354), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(G155gat), .B2(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(KEYINPUT77), .ZN(new_n374));
  XNOR2_X1  g173(.A(G141gat), .B(G148gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n376), .A2(KEYINPUT78), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n376), .A2(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT79), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G155gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n376), .B1(new_n384), .B2(G162gat), .ZN(new_n385));
  XOR2_X1   g184(.A(G141gat), .B(G148gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G155gat), .B(G162gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n374), .A2(new_n379), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n367), .B1(new_n268), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n263), .A2(new_n265), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n258), .A2(new_n255), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n257), .A2(new_n251), .A3(new_n253), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n392), .A2(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n381), .A2(new_n383), .ZN(new_n397));
  INV_X1    g196(.A(G162gat), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT2), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n373), .A2(new_n375), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n378), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n386), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n369), .B1(new_n387), .B2(new_n368), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n399), .A2(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(new_n404), .A3(KEYINPUT80), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n268), .A2(new_n389), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n366), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n393), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n389), .A2(KEYINPUT3), .B1(new_n410), .B2(new_n259), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n405), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n404), .A3(KEYINPUT4), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT4), .B1(new_n396), .B2(new_n404), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n390), .A2(new_n405), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT5), .B(new_n408), .C1(new_n411), .C2(new_n413), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n409), .A2(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  AOI21_X1  g226(.A(KEYINPUT6), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n418), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G228gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n331), .A2(new_n413), .B1(new_n316), .B2(new_n322), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n316), .A2(new_n331), .A3(new_n322), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n404), .B1(new_n441), .B2(new_n412), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g243(.A(KEYINPUT82), .B(new_n404), .C1(new_n441), .C2(new_n412), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n439), .B2(KEYINPUT81), .ZN(new_n447));
  INV_X1    g246(.A(new_n442), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n448), .C1(KEYINPUT81), .C2(new_n439), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT31), .B(G50gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n446), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n446), .B2(new_n449), .ZN(new_n453));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n446), .A2(new_n449), .A3(new_n451), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n365), .A2(new_n436), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n302), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n302), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n456), .B1(new_n452), .B2(new_n453), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n459), .A2(new_n455), .A3(new_n460), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n351), .B1(new_n363), .B2(KEYINPUT37), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n323), .B1(new_n355), .B2(new_n356), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT37), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n358), .A2(new_n323), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n434), .A2(new_n435), .A3(new_n359), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n363), .A2(KEYINPUT37), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT38), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n469), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n351), .B1(new_n342), .B2(new_n347), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n359), .A3(new_n361), .ZN(new_n483));
  OR4_X1    g282(.A1(new_n342), .A2(new_n347), .A3(new_n351), .A4(new_n353), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT84), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n411), .A2(new_n413), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n421), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n408), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n407), .A2(new_n408), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(KEYINPUT39), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT39), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n495), .A3(new_n408), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n427), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(KEYINPUT39), .A3(new_n493), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n496), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(new_n433), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n487), .A2(new_n488), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n464), .A2(new_n466), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n291), .A2(new_n292), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n505), .A2(new_n468), .A3(new_n467), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n365), .A2(KEYINPUT84), .ZN(new_n508));
  INV_X1    g307(.A(new_n488), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n434), .A2(new_n435), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n485), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n468), .A3(new_n467), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT35), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n504), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(KEYINPUT16), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n525));
  OAI21_X1  g324(.A(G8gat), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n522), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT88), .A3(G50gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n532), .B(new_n534), .C1(new_n536), .C2(KEYINPUT88), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT89), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT86), .Z(new_n542));
  NOR3_X1   g341(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT90), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n543), .B(KEYINPUT87), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n540), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT15), .A3(new_n535), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n531), .B1(new_n550), .B2(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n549), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n551), .A2(new_n554), .B1(new_n531), .B2(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT18), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  INV_X1    g357(.A(new_n554), .ZN(new_n559));
  INV_X1    g358(.A(new_n531), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n552), .B2(new_n553), .ZN(new_n561));
  OAI22_X1  g360(.A1(new_n559), .A2(new_n561), .B1(new_n560), .B2(new_n550), .ZN(new_n562));
  INV_X1    g361(.A(new_n556), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n560), .B(new_n552), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n556), .B(KEYINPUT13), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n557), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n557), .A2(new_n564), .A3(new_n575), .A4(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G57gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G64gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(G64gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(KEYINPUT94), .B2(new_n585), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(KEYINPUT94), .B2(new_n585), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n589), .A3(new_n583), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n560), .B1(new_n580), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT95), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n580), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G127gat), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n607), .A3(new_n608), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT41), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n614), .A2(new_n615), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT97), .B(G85gat), .Z(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT7), .ZN(new_n625));
  INV_X1    g424(.A(G99gat), .ZN(new_n626));
  INV_X1    g425(.A(G106gat), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT8), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G99gat), .B(G106gat), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n623), .A2(new_n632), .A3(new_n625), .A4(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n620), .B1(new_n552), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT98), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n550), .A2(KEYINPUT17), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n554), .A3(new_n634), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n639), .B1(new_n637), .B2(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n619), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n618), .A3(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT99), .B1(new_n595), .B2(new_n634), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n591), .A2(new_n631), .A3(new_n594), .A4(new_n633), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n635), .A2(KEYINPUT99), .A3(new_n591), .A4(new_n594), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n649), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G120gat), .B(G148gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT100), .ZN(new_n661));
  XOR2_X1   g460(.A(G176gat), .B(G204gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n612), .A2(new_n648), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n436), .A2(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n436), .A2(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n516), .A2(new_n579), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  AOI22_X1  g474(.A1(new_n463), .A2(KEYINPUT83), .B1(new_n481), .B2(new_n502), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n676), .A2(new_n466), .B1(new_n514), .B2(new_n510), .ZN(new_n677));
  INV_X1    g476(.A(new_n579), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n508), .A2(new_n509), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n677), .A2(new_n678), .A3(new_n680), .A4(new_n668), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n528), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  NOR3_X1   g485(.A1(new_n677), .A2(new_n678), .A3(new_n668), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n687), .B2(new_n505), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n301), .A2(G15gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT102), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n687), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n469), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n648), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n612), .A2(new_n678), .A3(new_n666), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G29gat), .A3(new_n672), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n677), .B2(new_n648), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n481), .A2(new_n502), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n457), .A2(new_n461), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n483), .A2(new_n484), .B1(new_n435), .B2(new_n434), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT105), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n512), .A2(new_n707), .A3(new_n469), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n302), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n515), .B1(new_n703), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n645), .A2(new_n647), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n712));
  AND4_X1   g511(.A1(new_n702), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n301), .B1(new_n462), .B2(KEYINPUT105), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n503), .A2(new_n714), .A3(new_n708), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n648), .B1(new_n715), .B2(new_n515), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n702), .B1(new_n716), .B2(new_n712), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n701), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n697), .B(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n672), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n700), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n698), .A2(G36gat), .A3(new_n680), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n680), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n720), .B2(new_n302), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n696), .A2(new_n533), .A3(new_n505), .A4(new_n697), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(KEYINPUT47), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1330gat));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n698), .A2(G50gat), .A3(new_n704), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n469), .A3(new_n719), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  INV_X1    g540(.A(new_n719), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n702), .A3(new_n712), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n742), .B1(new_n746), .B2(new_n701), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n741), .B1(new_n747), .B2(new_n469), .ZN(new_n748));
  OAI211_X1 g547(.A(KEYINPUT108), .B(new_n734), .C1(new_n748), .C2(new_n736), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n740), .A2(new_n749), .ZN(G1331gat));
  NAND4_X1  g549(.A1(new_n612), .A2(new_n678), .A3(new_n648), .A4(new_n666), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n515), .B2(new_n715), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n671), .B(KEYINPUT110), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g555(.A1(new_n752), .A2(new_n679), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT111), .ZN(G1333gat));
  NAND2_X1  g561(.A1(new_n752), .A2(new_n301), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n291), .A2(new_n292), .A3(G71gat), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n763), .A2(G71gat), .B1(new_n752), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n752), .A2(new_n469), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n612), .A2(new_n579), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n711), .A4(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n710), .A2(new_n711), .A3(new_n769), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n776), .A2(new_n621), .A3(new_n666), .A4(new_n671), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n516), .A2(new_n711), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n744), .A2(new_n745), .B1(new_n778), .B2(KEYINPUT44), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n769), .A2(new_n666), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n672), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n783), .B2(new_n621), .ZN(G1336gat));
  NOR3_X1   g583(.A1(new_n779), .A2(new_n680), .A3(new_n780), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n680), .A2(G92gat), .A3(new_n667), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT51), .B1(new_n773), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n788), .B2(new_n773), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n772), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n786), .A2(G92gat), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n770), .A2(new_n771), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n771), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n795), .A2(new_n796), .B1(new_n774), .B2(new_n773), .ZN(new_n797));
  INV_X1    g596(.A(new_n787), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n776), .A2(KEYINPUT114), .A3(new_n787), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n793), .B1(new_n785), .B2(new_n622), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n792), .A2(new_n793), .B1(new_n801), .B2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n782), .B2(new_n302), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n666), .A2(new_n626), .A3(new_n505), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n797), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n704), .A2(new_n667), .A3(G106gat), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n791), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n627), .B1(new_n781), .B2(new_n469), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n776), .A2(new_n807), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n811), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n810), .A2(new_n811), .B1(new_n813), .B2(new_n809), .ZN(G1339gat));
  NAND4_X1  g613(.A1(new_n612), .A2(new_n678), .A3(new_n648), .A4(new_n667), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n555), .B2(new_n556), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n565), .A2(KEYINPUT116), .A3(new_n567), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n565), .A2(new_n567), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n555), .A2(new_n817), .A3(new_n556), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n573), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n578), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n649), .C1(new_n654), .C2(new_n656), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n663), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n658), .A2(new_n655), .ZN(new_n831));
  INV_X1    g630(.A(new_n656), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(G230gat), .A3(G233gat), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n834), .A3(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n664), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n830), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n826), .A2(new_n711), .A3(new_n827), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n825), .A2(new_n647), .A3(new_n645), .A4(new_n578), .ZN(new_n840));
  INV_X1    g639(.A(new_n838), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n579), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n578), .A3(new_n666), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n839), .B(new_n842), .C1(new_n845), .C2(new_n711), .ZN(new_n846));
  INV_X1    g645(.A(new_n612), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n816), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n848), .A2(new_n513), .A3(new_n679), .A4(new_n753), .ZN(new_n849));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n579), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n839), .A2(new_n842), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n711), .B1(new_n843), .B2(new_n844), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n815), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n704), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n848), .B2(new_n469), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n672), .A2(new_n679), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n505), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n678), .A2(new_n255), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(G1340gat));
  INV_X1    g662(.A(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(G120gat), .B1(new_n864), .B2(new_n667), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n666), .A2(new_n258), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT119), .Z(new_n867));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n864), .B2(new_n847), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n849), .A2(new_n252), .A3(new_n612), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n864), .B2(new_n648), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n849), .A2(new_n250), .A3(new_n711), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n302), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT120), .Z(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n854), .B2(new_n469), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n469), .A2(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n836), .B2(new_n837), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n830), .A2(new_n834), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n664), .A4(new_n835), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n579), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n711), .B1(new_n888), .B2(new_n844), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n847), .B1(new_n851), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n881), .B1(new_n890), .B2(new_n815), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n579), .B(new_n878), .C1(new_n879), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n302), .A2(new_n469), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n848), .A2(new_n679), .A3(new_n753), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n678), .A2(G141gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n893), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n895), .B1(new_n893), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n840), .A2(new_n841), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n847), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n815), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n704), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n815), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n848), .A2(new_n881), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n878), .A2(new_n666), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT59), .B(G148gat), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n914), .A3(new_n666), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n879), .A2(new_n891), .ZN(new_n916));
  INV_X1    g715(.A(new_n878), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n918), .B2(new_n666), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n913), .B(new_n915), .C1(new_n919), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n397), .A3(new_n612), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n916), .A2(new_n847), .A3(new_n917), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n397), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n897), .B2(new_n711), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n648), .A2(new_n398), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n918), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n848), .A2(new_n671), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n680), .A2(new_n513), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n929), .A2(new_n579), .A3(new_n235), .A4(new_n236), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n753), .A2(new_n505), .A3(new_n679), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n856), .B2(new_n857), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n579), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n206), .ZN(G1348gat));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n207), .A3(new_n666), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n932), .A2(new_n666), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n207), .ZN(G1349gat));
  AOI21_X1  g736(.A(new_n219), .B1(new_n932), .B2(new_n612), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n929), .A2(new_n215), .A3(new_n612), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT124), .B(KEYINPUT60), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n929), .A2(new_n215), .A3(new_n612), .ZN(new_n941));
  NAND2_X1  g740(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n932), .A2(new_n612), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(new_n219), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n940), .A2(new_n944), .ZN(G1350gat));
  AOI211_X1 g744(.A(new_n648), .B(new_n931), .C1(new_n856), .C2(new_n857), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n946), .A2(new_n947), .A3(new_n217), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(new_n217), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n927), .A2(new_n217), .A3(new_n711), .A4(new_n928), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT125), .Z(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n680), .A2(new_n896), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT126), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n927), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n579), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n753), .A2(new_n679), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n911), .A2(new_n301), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n579), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  OR2_X1    g759(.A1(new_n909), .A2(new_n910), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n957), .A2(new_n301), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n666), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n667), .A2(G204gat), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n955), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n955), .A2(new_n966), .ZN(new_n968));
  XNOR2_X1  g767(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n964), .A2(new_n970), .ZN(G1353gat));
  INV_X1    g770(.A(new_n955), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n972), .A2(new_n317), .A3(new_n847), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n612), .B(new_n962), .C1(new_n909), .C2(new_n910), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n711), .A3(new_n962), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G218gat), .ZN(new_n979));
  OR3_X1    g778(.A1(new_n972), .A2(G218gat), .A3(new_n648), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1355gat));
endmodule


