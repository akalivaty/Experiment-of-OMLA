//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n218), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n222), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OAI22_X1  g0047(.A1(new_n247), .A2(new_n209), .B1(new_n223), .B2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n223), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(new_n202), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n245), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT11), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n252), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n245), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G68), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n253), .A2(new_n254), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(G274), .B1(new_n269), .B2(new_n222), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n275), .B2(G238), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n279), .A2(new_n283), .A3(G226), .A4(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n279), .A2(new_n283), .A3(G232), .A4(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  INV_X1    g0089(.A(new_n273), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n276), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n276), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(G169), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(G179), .A3(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n297), .B2(G169), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n264), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n279), .A2(new_n283), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G222), .A3(new_n284), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G223), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n305), .B1(new_n202), .B2(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n290), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n271), .B1(new_n275), .B2(G226), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n223), .B1(new_n201), .B2(new_n203), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n315), .A2(new_n249), .B1(new_n316), .B2(new_n247), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n245), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n261), .A2(G50), .A3(new_n262), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(G50), .C2(new_n256), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT9), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n309), .A2(G190), .A3(new_n310), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT70), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT10), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n321), .A2(new_n323), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT10), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n322), .A3(new_n327), .A4(new_n312), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n315), .B1(KEYINPUT69), .B2(new_n247), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(KEYINPUT69), .B2(new_n247), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n331), .B1(new_n223), .B2(new_n202), .C1(new_n249), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n245), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n202), .B1(new_n255), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n261), .A2(new_n335), .B1(new_n202), .B2(new_n257), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G274), .ZN(new_n338));
  AND2_X1   g0138(.A1(G1), .A2(G13), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n272), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n267), .ZN(new_n341));
  INV_X1    g0141(.A(G244), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n274), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n304), .A2(G232), .A3(new_n284), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  INV_X1    g0145(.A(G238), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n344), .B1(new_n345), .B2(new_n304), .C1(new_n306), .C2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n347), .B2(new_n290), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n337), .B1(new_n348), .B2(G169), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n337), .B1(new_n348), .B2(G190), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n329), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n311), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n320), .C1(G179), .C2(new_n311), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT68), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n264), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n297), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n355), .B1(new_n294), .B2(new_n296), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n261), .ZN(new_n370));
  INV_X1    g0170(.A(new_n315), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n262), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n370), .A2(new_n372), .B1(new_n256), .B2(new_n371), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n277), .A2(new_n278), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n210), .A2(G1698), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(G223), .C2(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n273), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n341), .B1(new_n274), .B2(new_n229), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n355), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n290), .ZN(new_n383));
  INV_X1    g0183(.A(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(G190), .ZN(new_n386));
  INV_X1    g0186(.A(G58), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n258), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n203), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n246), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n281), .A2(new_n282), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n279), .B2(new_n283), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(KEYINPUT7), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(G68), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n375), .B2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n393), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n391), .B1(new_n400), .B2(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n245), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n374), .B(new_n386), .C1(new_n397), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n245), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(KEYINPUT16), .B2(new_n396), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n374), .A4(new_n386), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n406), .A2(KEYINPUT72), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT72), .B1(new_n406), .B2(new_n410), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  INV_X1    g0213(.A(new_n393), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n279), .A2(new_n283), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n223), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n398), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n258), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n373), .B1(new_n420), .B2(new_n408), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n379), .A2(new_n380), .A3(new_n351), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G169), .B2(new_n385), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n409), .A2(new_n374), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  INV_X1    g0226(.A(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n411), .A2(new_n412), .A3(new_n429), .ZN(new_n430));
  AND4_X1   g0230(.A1(new_n303), .A2(new_n363), .A3(new_n369), .A4(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n284), .B1(new_n277), .B2(new_n278), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n415), .A2(G303), .B1(G264), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT80), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n375), .A2(new_n434), .A3(G257), .A4(new_n284), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n284), .A2(G257), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT80), .B1(new_n392), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n290), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n266), .A2(G1), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n446), .B2(new_n270), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n255), .A2(G45), .ZN(new_n448));
  OR2_X1    g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(KEYINPUT73), .A3(new_n340), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n446), .A2(G270), .A3(new_n273), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT21), .A3(G169), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n440), .B(G179), .C1(new_n455), .C2(new_n456), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n245), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(G33), .B2(G283), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(G33), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n466), .A2(KEYINPUT82), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n464), .B2(new_n465), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n467), .A2(KEYINPUT82), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n467), .A2(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n256), .A2(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n255), .A2(G33), .ZN(new_n477));
  AND4_X1   g0277(.A1(new_n222), .A2(new_n256), .A3(new_n244), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(G116), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n471), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n460), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n480), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n458), .B2(new_n459), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n446), .A2(new_n270), .A3(new_n441), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT73), .B1(new_n450), .B2(new_n340), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n454), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT79), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n359), .B1(new_n492), .B2(new_n440), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n480), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n273), .B1(new_n433), .B2(new_n438), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n490), .B2(new_n491), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G190), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n484), .B(new_n499), .C1(new_n355), .C2(new_n498), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n483), .A2(new_n486), .A3(new_n496), .A4(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n446), .A2(G264), .A3(new_n273), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n284), .C1(new_n281), .C2(new_n282), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n432), .A2(KEYINPUT87), .A3(G257), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n452), .B(new_n503), .C1(new_n511), .C2(new_n273), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n359), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n504), .A2(new_n505), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT87), .B1(new_n432), .B2(G257), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n508), .A2(new_n509), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n290), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n351), .A3(new_n452), .A4(new_n503), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n211), .A2(KEYINPUT22), .A3(G20), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n279), .A2(new_n283), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n279), .A2(new_n283), .A3(new_n524), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n375), .A2(new_n223), .A3(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n223), .B1(new_n531), .B2(KEYINPUT23), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n345), .A3(G20), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(KEYINPUT85), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n533), .B2(new_n345), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(KEYINPUT24), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n523), .A2(new_n525), .B1(KEYINPUT22), .B2(new_n527), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n543), .A3(new_n245), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n257), .A2(new_n345), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT86), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT25), .ZN(new_n547));
  XOR2_X1   g0347(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n548));
  INV_X1    g0348(.A(new_n478), .ZN(new_n549));
  OAI221_X1 g0349(.A(new_n547), .B1(new_n545), .B2(new_n548), .C1(new_n549), .C2(new_n345), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n520), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n529), .A2(new_n538), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n407), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n554), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n512), .A2(new_n355), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G190), .B2(new_n512), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n552), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n346), .A2(new_n284), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n342), .A2(G1698), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n281), .C2(new_n282), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n273), .B1(new_n561), .B2(new_n530), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n273), .A2(G274), .A3(new_n442), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n212), .B1(new_n255), .B2(G45), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n273), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT77), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n340), .A2(new_n442), .B1(new_n273), .B2(new_n564), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT77), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G238), .A2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n342), .B2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n531), .B1(new_n571), .B2(new_n375), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n568), .B(new_n569), .C1(new_n572), .C2(new_n273), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(new_n573), .A3(G200), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n223), .B1(new_n287), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(G97), .A2(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n211), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n223), .B(G68), .C1(new_n281), .C2(new_n282), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n575), .B1(new_n249), .B2(new_n469), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n245), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n332), .A2(new_n257), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n478), .A2(G87), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n567), .A2(new_n573), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(KEYINPUT78), .B1(G190), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT78), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n574), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n351), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n583), .B(new_n584), .C1(new_n332), .C2(new_n549), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n567), .A2(new_n573), .A3(new_n359), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n589), .A2(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n558), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(new_n284), .C1(new_n281), .C2(new_n282), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(G33), .B2(G283), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n279), .A2(new_n283), .A3(G250), .A4(G1698), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n342), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n279), .A2(new_n283), .A3(new_n284), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n290), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n450), .A2(new_n290), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n447), .A2(new_n451), .B1(new_n606), .B2(G257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n359), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n256), .A2(G97), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n478), .B2(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n246), .A2(G77), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n613), .A2(new_n469), .A3(G107), .ZN(new_n614));
  XNOR2_X1  g0414(.A(G97), .B(G107), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n616), .B2(new_n223), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n395), .B2(G107), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n611), .B1(new_n618), .B2(new_n407), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n605), .A2(new_n351), .A3(new_n607), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n609), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT76), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT76), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n609), .A2(new_n619), .A3(new_n623), .A4(new_n620), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n605), .A2(G190), .A3(new_n607), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT74), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT74), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n605), .A2(new_n627), .A3(G190), .A4(new_n607), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n355), .B1(new_n605), .B2(new_n607), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT75), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n629), .B2(new_n631), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n622), .B(new_n624), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n501), .A2(new_n597), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n431), .A2(new_n636), .ZN(G372));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  INV_X1    g0438(.A(new_n621), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n561), .A2(new_n530), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n290), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT88), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n563), .A2(new_n565), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n563), .B2(new_n565), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n359), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n592), .A2(new_n593), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n569), .B1(new_n641), .B2(new_n568), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n562), .A2(new_n566), .A3(KEYINPUT77), .ZN(new_n649));
  OAI21_X1  g0449(.A(G190), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(G200), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n586), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n647), .B2(new_n652), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n638), .B(new_n639), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n647), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n622), .A2(new_n624), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n638), .B1(new_n658), .B2(new_n596), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n552), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n481), .A3(new_n496), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n629), .A2(new_n631), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT75), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n647), .A2(new_n652), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n555), .B2(new_n557), .ZN(new_n670));
  INV_X1    g0470(.A(new_n658), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n662), .A2(new_n666), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n431), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n429), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n349), .B1(new_n351), .B2(new_n348), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n297), .A2(G169), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT14), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n300), .A3(new_n299), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n369), .A2(new_n676), .B1(new_n679), .B2(new_n264), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n411), .A2(new_n412), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n675), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n362), .B1(new_n683), .B2(new_n329), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n674), .A2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n255), .A2(new_n223), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n496), .B1(new_n485), .B2(KEYINPUT83), .ZN(new_n692));
  AOI211_X1 g0492(.A(new_n482), .B(new_n484), .C1(new_n458), .C2(new_n459), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n558), .B1(new_n555), .B2(new_n691), .ZN(new_n695));
  INV_X1    g0495(.A(new_n691), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n552), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT91), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT91), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n694), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n661), .A2(new_n696), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n484), .A2(new_n691), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT21), .B1(new_n493), .B2(new_n480), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n485), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n501), .B2(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n219), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n577), .A2(new_n211), .A3(new_n461), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n255), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n226), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n483), .A2(new_n486), .A3(new_n496), .A4(new_n661), .ZN(new_n720));
  INV_X1    g0520(.A(new_n635), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n670), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n639), .B1(new_n654), .B2(new_n655), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT26), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n658), .A2(new_n638), .A3(new_n596), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n724), .A2(new_n647), .A3(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n719), .B(new_n696), .C1(new_n722), .C2(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n723), .A2(KEYINPUT26), .B1(new_n594), .B2(new_n646), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n692), .A2(new_n693), .A3(new_n552), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n666), .A2(new_n670), .A3(new_n671), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n725), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT94), .B1(new_n731), .B2(new_n691), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT29), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n696), .B1(new_n660), .B2(new_n672), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n500), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n692), .A2(new_n693), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n558), .A2(new_n596), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n721), .A4(new_n691), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n645), .A2(new_n351), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n457), .A2(new_n608), .A3(new_n512), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n588), .A2(new_n518), .A3(new_n503), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n605), .A2(new_n607), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n498), .A3(G179), .A4(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT92), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n502), .B1(new_n517), .B2(new_n290), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n605), .A3(new_n588), .A4(new_n607), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n459), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT92), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n743), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n747), .B1(new_n459), .B2(new_n750), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n691), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n752), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n459), .A2(new_n750), .A3(KEYINPUT92), .A4(new_n747), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n742), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n746), .A2(new_n763), .A3(new_n747), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(KEYINPUT93), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n696), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n757), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n740), .A2(new_n759), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G330), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n736), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n718), .B1(new_n772), .B2(G1), .ZN(G364));
  INV_X1    g0573(.A(G13), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n255), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n714), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n710), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n708), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n222), .B1(G20), .B2(new_n359), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n223), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n365), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G107), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n304), .C1(new_n211), .C2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT96), .Z(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT32), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n223), .A2(new_n351), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(new_n365), .A3(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n790), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(new_n258), .B2(new_n797), .C1(new_n202), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(G190), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n387), .B1(new_n794), .B2(new_n793), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n365), .A2(G179), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n223), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n800), .A2(new_n355), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n809), .B2(new_n209), .ZN(new_n810));
  OR4_X1    g0610(.A1(new_n789), .A2(new_n799), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n798), .ZN(new_n812));
  INV_X1    g0612(.A(new_n791), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n812), .B1(new_n813), .B2(G329), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT33), .B(G317), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n797), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G294), .A2(new_n806), .B1(new_n801), .B2(G322), .ZN(new_n818));
  INV_X1    g0618(.A(new_n787), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n808), .A2(G326), .B1(new_n819), .B2(G303), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n304), .B1(G283), .B2(new_n785), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n782), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n781), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n239), .A2(G45), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n713), .A2(new_n375), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n266), .B2(new_n226), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n713), .A2(new_n415), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G355), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(G116), .B2(new_n219), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT95), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n829), .A2(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n778), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n823), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n826), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n708), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n780), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  NAND3_X1  g0645(.A1(new_n350), .A2(new_n352), .A3(new_n691), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n354), .A2(new_n356), .B1(new_n337), .B2(new_n696), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n676), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n734), .B(new_n849), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n850), .A2(new_n770), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n778), .B1(new_n850), .B2(new_n770), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n782), .A2(new_n825), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n778), .B1(G77), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n849), .A2(new_n825), .ZN(new_n856));
  INV_X1    g0656(.A(G294), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n802), .A2(new_n857), .B1(new_n345), .B2(new_n787), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G116), .A2(new_n812), .B1(new_n813), .B2(G311), .ZN(new_n859));
  XOR2_X1   g0659(.A(KEYINPUT97), .B(G283), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n797), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(G303), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n809), .A2(new_n862), .B1(new_n211), .B2(new_n784), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n807), .A2(new_n415), .ZN(new_n864));
  OR4_X1    g0664(.A1(new_n858), .A2(new_n861), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n375), .B1(new_n791), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G68), .B2(new_n785), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n806), .A2(G58), .B1(new_n819), .B2(G50), .ZN(new_n869));
  INV_X1    g0669(.A(new_n797), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(G150), .B1(new_n812), .B2(G159), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT98), .B(G143), .Z(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(new_n802), .B2(new_n872), .C1(new_n873), .C2(new_n809), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT34), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n868), .B(new_n869), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n865), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n855), .B(new_n856), .C1(new_n781), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n853), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n775), .A2(new_n255), .ZN(new_n882));
  INV_X1    g0682(.A(new_n689), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n429), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n374), .B1(new_n403), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n427), .B2(new_n689), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n404), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n425), .A2(new_n427), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n425), .A2(new_n689), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n404), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n886), .A2(new_n689), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n430), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT38), .B(new_n894), .C1(new_n430), .C2(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n485), .A2(new_n552), .A3(new_n706), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n557), .A2(new_n544), .A3(new_n551), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n654), .B2(new_n655), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n635), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n591), .A3(new_n650), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n592), .A2(new_n595), .A3(new_n593), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n622), .B2(new_n624), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n647), .B(new_n656), .C1(new_n909), .C2(new_n638), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n691), .B(new_n849), .C1(new_n904), .C2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n846), .B(KEYINPUT99), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n691), .A2(new_n364), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n679), .B2(new_n368), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(KEYINPUT100), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n303), .A2(new_n369), .A3(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n911), .A2(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n900), .B1(new_n918), .B2(KEYINPUT101), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n915), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n696), .B(new_n848), .C1(new_n660), .C2(new_n672), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT101), .B(new_n920), .C1(new_n921), .C2(new_n912), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n884), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT102), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT101), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n912), .B1(new_n734), .B2(new_n849), .ZN(new_n927));
  INV_X1    g0727(.A(new_n920), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n922), .A3(new_n900), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT102), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(new_n884), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n679), .A2(new_n264), .A3(new_n691), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n404), .B1(new_n421), .B2(new_n423), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n421), .A2(new_n883), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(KEYINPUT103), .A3(new_n893), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT103), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(KEYINPUT37), .C1(new_n934), .C2(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n406), .A2(new_n410), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n935), .B1(new_n429), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n897), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT104), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n899), .A3(new_n898), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n899), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n944), .A2(KEYINPUT39), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n933), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n925), .A2(new_n932), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n733), .A2(new_n431), .A3(new_n735), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n684), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n848), .B1(new_n917), .B2(new_n915), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n755), .B(new_n763), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n691), .B1(new_n754), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT31), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT105), .B1(new_n767), .B2(new_n757), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n754), .A2(new_n959), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n758), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n740), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n948), .B(new_n958), .C1(new_n964), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT40), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT40), .B1(new_n898), .B2(new_n899), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n740), .A2(new_n966), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n961), .B1(new_n960), .B2(KEYINPUT31), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n767), .A2(KEYINPUT105), .A3(new_n757), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(new_n975), .A3(new_n958), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n431), .A2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  INV_X1    g0781(.A(G330), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n882), .B1(new_n957), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n957), .B2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(new_n616), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT35), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT35), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n988), .A2(G116), .A3(new_n224), .A4(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT36), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n226), .B(G77), .C1(new_n387), .C2(new_n258), .ZN(new_n992));
  INV_X1    g0792(.A(new_n201), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n258), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(G1), .A3(new_n774), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n986), .A2(new_n991), .A3(new_n995), .ZN(G367));
  OR2_X1    g0796(.A1(new_n691), .A2(new_n586), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n647), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n668), .A2(new_n669), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n696), .A2(new_n619), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n721), .A2(new_n1001), .B1(new_n639), .B2(new_n696), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT42), .B1(new_n701), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n701), .A2(KEYINPUT42), .A3(new_n1003), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n671), .B1(new_n1002), .B2(new_n661), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1005), .A2(new_n1006), .B1(new_n691), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1000), .B1(new_n1008), .B2(KEYINPUT106), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n691), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1006), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n1004), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT106), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1000), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1009), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT43), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n711), .A2(new_n1002), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n1016), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n1025), .B2(new_n1018), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n703), .B2(new_n1003), .ZN(new_n1029));
  OAI211_X1 g0829(.A(KEYINPUT44), .B(new_n1002), .C1(new_n701), .C2(new_n702), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n694), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n704), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n702), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n1003), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n711), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT108), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1031), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1044), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1039), .A2(new_n1031), .A3(new_n1046), .A4(new_n1042), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1033), .A2(KEYINPUT107), .A3(new_n709), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT107), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n710), .B1(new_n701), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n704), .A2(new_n1032), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n771), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n771), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n714), .B(KEYINPUT41), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n776), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1027), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(G317), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n392), .B1(new_n791), .B2(new_n1060), .C1(new_n469), .C2(new_n784), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT109), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n860), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G294), .A2(new_n870), .B1(new_n1063), .B2(new_n812), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n345), .B2(new_n805), .ZN(new_n1065));
  INV_X1    g0865(.A(G311), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n802), .A2(new_n862), .B1(new_n809), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n787), .A2(new_n461), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT46), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1062), .A2(new_n1065), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT110), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G68), .A2(new_n806), .B1(new_n801), .B2(G150), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT111), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n797), .A2(new_n792), .B1(new_n791), .B2(new_n873), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n993), .B2(new_n812), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n415), .B1(G77), .B2(new_n785), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n872), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n808), .A2(new_n1077), .B1(new_n819), .B2(G58), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1071), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT47), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n781), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n827), .B1(new_n219), .B2(new_n332), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n830), .B2(new_n235), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n840), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(new_n842), .C2(new_n1014), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1059), .A2(new_n1086), .ZN(G387));
  INV_X1    g0887(.A(new_n1054), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n699), .A2(new_n700), .A3(new_n826), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n798), .A2(new_n258), .B1(new_n791), .B2(new_n316), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n392), .B(new_n1090), .C1(new_n371), .C2(new_n870), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n787), .A2(new_n202), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n805), .A2(new_n332), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G50), .C2(new_n801), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n808), .A2(G159), .B1(new_n785), .B2(G97), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n375), .B1(new_n813), .B2(G326), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n805), .A2(new_n860), .B1(new_n787), .B2(new_n857), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n870), .A2(G311), .B1(new_n812), .B2(G303), .ZN(new_n1099));
  INV_X1    g0899(.A(G322), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1099), .B1(new_n802), .B2(new_n1060), .C1(new_n1100), .C2(new_n809), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT49), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1097), .B1(new_n461), .B2(new_n784), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1096), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT112), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n782), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n232), .A2(new_n266), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n830), .B1(new_n715), .B2(new_n833), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT50), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n371), .B2(new_n209), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n315), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n266), .B1(new_n258), .B2(new_n202), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n715), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1113), .A2(new_n1118), .B1(G107), .B2(new_n219), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n840), .B1(new_n1119), .B2(new_n827), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1111), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT113), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1088), .A2(new_n777), .B1(new_n1089), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1088), .A2(new_n772), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n714), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1088), .A2(new_n772), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(G393));
  INV_X1    g0927(.A(KEYINPUT118), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1124), .A2(new_n1045), .A3(KEYINPUT118), .A4(new_n1047), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n714), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1048), .A2(new_n777), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n827), .B1(new_n469), .B2(new_n219), .C1(new_n831), .C2(new_n242), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n778), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G150), .A2(new_n808), .B1(new_n801), .B2(G159), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT51), .Z(new_n1141));
  AOI22_X1  g0941(.A1(new_n870), .A2(new_n993), .B1(new_n812), .B2(new_n371), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n806), .A2(G77), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n392), .B1(new_n1077), .B2(new_n813), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n258), .B2(new_n787), .C1(new_n211), .C2(new_n784), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT115), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G311), .A2(new_n801), .B1(new_n808), .B2(G317), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT52), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n798), .A2(new_n857), .B1(new_n791), .B2(new_n1100), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G303), .B2(new_n870), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n806), .A2(G116), .B1(new_n1063), .B2(new_n819), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1153), .A2(new_n415), .A3(new_n786), .A4(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1146), .A2(new_n1149), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1137), .B(new_n1139), .C1(new_n781), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1003), .B2(new_n842), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1134), .A2(new_n1135), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n776), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1158), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT117), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1131), .A2(new_n1133), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G390));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n933), .B1(new_n927), .B2(new_n928), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n947), .A2(new_n951), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n769), .A2(G330), .A3(new_n920), .A4(new_n849), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n847), .A2(new_n676), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n727), .B2(new_n732), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n928), .B1(new_n1171), .B2(new_n846), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n948), .A2(new_n933), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1167), .B(new_n1168), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n724), .A2(new_n647), .A3(new_n725), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n730), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n720), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n719), .B1(new_n1177), .B2(new_n696), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n731), .A2(KEYINPUT94), .A3(new_n691), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1169), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n846), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n920), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1173), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n950), .B1(KEYINPUT39), .B2(new_n946), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1182), .A2(new_n1183), .B1(new_n1184), .B2(new_n1166), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n982), .B1(new_n971), .B2(new_n974), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n958), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1174), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n431), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n955), .A2(new_n684), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1171), .A2(new_n846), .A3(new_n1168), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n920), .B1(new_n1186), .B2(new_n849), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n769), .A2(G330), .A3(new_n849), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1186), .A2(new_n958), .B1(new_n1194), .B2(new_n928), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1192), .A2(new_n1193), .B1(new_n1195), .B2(new_n927), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1165), .B1(new_n1188), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1186), .A2(new_n849), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1168), .C1(new_n1200), .C2(new_n920), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1194), .A2(new_n928), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1187), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n927), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1190), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1167), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n958), .A3(new_n1186), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1208), .A3(KEYINPUT119), .A4(new_n1174), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1198), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1197), .A2(KEYINPUT120), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1188), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n714), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT121), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1188), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1184), .A2(new_n824), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n778), .B1(new_n371), .B2(new_n854), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n797), .A2(new_n345), .B1(new_n798), .B2(new_n469), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G294), .B2(new_n813), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n304), .B1(G87), .B2(new_n819), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n806), .A2(G77), .B1(new_n785), .B2(G68), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G116), .A2(new_n801), .B1(new_n808), .B2(G283), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n802), .A2(new_n866), .B1(new_n201), .B2(new_n784), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G159), .B2(new_n806), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n813), .A2(G125), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT54), .B(G143), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n870), .A2(G137), .B1(new_n812), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n415), .B1(new_n808), .B2(G128), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1227), .A2(new_n1228), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n819), .A2(G150), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT53), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1225), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1219), .B1(new_n1236), .B2(new_n781), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1217), .A2(new_n777), .B1(new_n1218), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1215), .A2(new_n1216), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1216), .B1(new_n1215), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(G378));
  NAND2_X1  g1041(.A1(new_n1210), .A2(new_n1191), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n925), .A2(KEYINPUT123), .A3(new_n932), .A4(new_n953), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n329), .A2(new_n361), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n320), .A3(new_n689), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n320), .A2(new_n689), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n329), .A2(new_n361), .A3(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n920), .A2(new_n849), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n974), .B2(new_n971), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1253), .A2(new_n970), .B1(new_n968), .B2(KEYINPUT40), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1254), .B2(new_n982), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n977), .A2(G330), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1243), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n952), .B1(new_n924), .B2(KEYINPUT102), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT123), .B1(new_n1260), .B2(new_n932), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n930), .A2(new_n931), .A3(new_n884), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n931), .B1(new_n930), .B2(new_n884), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n952), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1265), .A2(new_n1258), .A3(KEYINPUT123), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1242), .A2(new_n1267), .A3(KEYINPUT57), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT57), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1190), .B1(new_n1198), .B2(new_n1209), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT122), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1256), .B1(new_n977), .B2(G330), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n982), .B(new_n1251), .C1(new_n969), .C2(new_n976), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1265), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1258), .A2(new_n954), .A3(new_n1271), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1268), .A2(new_n714), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1251), .A2(new_n824), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n778), .B1(new_n993), .B2(new_n854), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n797), .A2(new_n866), .B1(new_n798), .B2(new_n873), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G150), .A2(new_n806), .B1(new_n808), .B2(G125), .ZN(new_n1283));
  INV_X1    g1083(.A(G128), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n802), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1282), .B(new_n1285), .C1(new_n819), .C2(new_n1230), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT59), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n785), .A2(G159), .ZN(new_n1290));
  AOI211_X1 g1090(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n392), .B2(new_n265), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n802), .A2(new_n345), .B1(new_n387), .B2(new_n784), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G116), .B2(new_n808), .ZN(new_n1296));
  AOI211_X1 g1096(.A(G41), .B(new_n375), .C1(new_n870), .C2(G97), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n332), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1298), .A2(new_n812), .B1(new_n813), .B2(G283), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1092), .B1(G68), .B2(new_n806), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT58), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1292), .B(new_n1303), .C1(new_n1302), .C2(new_n1301), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1281), .B1(new_n1304), .B2(new_n781), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1280), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1277), .B2(new_n776), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1279), .A2(new_n1308), .ZN(G375));
  NOR2_X1   g1109(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1057), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1212), .A2(new_n1311), .A3(new_n1213), .A4(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n928), .A2(new_n824), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n778), .B1(G68), .B2(new_n854), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n797), .A2(new_n461), .B1(new_n791), .B2(new_n862), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(G107), .B2(new_n812), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1093), .B1(G283), .B2(new_n801), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n304), .B1(G77), .B2(new_n785), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n808), .A2(G294), .B1(new_n819), .B2(G97), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .A4(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(G132), .A2(new_n808), .B1(new_n801), .B2(G137), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n870), .A2(new_n1230), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n392), .B1(new_n812), .B2(G150), .ZN(new_n1324));
  AOI22_X1  g1124(.A1(new_n806), .A2(G50), .B1(new_n785), .B2(G58), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  OAI22_X1  g1126(.A1(new_n787), .A2(new_n792), .B1(new_n791), .B2(new_n1284), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(KEYINPUT124), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1321), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1315), .B1(new_n1329), .B2(new_n781), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1196), .A2(new_n777), .B1(new_n1314), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1313), .A2(new_n1331), .ZN(G381));
  OR2_X1    g1132(.A1(G393), .A2(G396), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1215), .A2(new_n1238), .ZN(new_n1334));
  NOR4_X1   g1134(.A1(new_n1333), .A2(new_n1334), .A3(G384), .A4(G381), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1086), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1269), .B1(new_n1210), .B2(new_n1191), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1132), .B1(new_n1338), .B2(new_n1267), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1307), .B1(new_n1339), .B2(new_n1278), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1335), .A2(new_n1337), .A3(new_n1340), .A4(new_n1163), .ZN(G407));
  INV_X1    g1141(.A(new_n1334), .ZN(new_n1342));
  INV_X1    g1142(.A(G343), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(G213), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1340), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(G407), .A2(G213), .A3(new_n1346), .ZN(G409));
  XNOR2_X1  g1147(.A(G393), .B(new_n844), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1348), .B1(G387), .B2(G390), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1337), .A2(new_n1163), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT126), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(G393), .B(G396), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1352), .B1(new_n1337), .B2(new_n1163), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1350), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT126), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G387), .A2(KEYINPUT127), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1348), .B1(new_n1357), .B2(G390), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(G387), .A2(KEYINPUT127), .A3(new_n1163), .ZN(new_n1359));
  AOI22_X1  g1159(.A1(new_n1351), .A2(new_n1356), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1132), .B1(new_n1310), .B2(KEYINPUT60), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT60), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1206), .A2(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(KEYINPUT125), .B1(new_n1364), .B2(new_n1310), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1197), .A2(KEYINPUT60), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT125), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1311), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1362), .B1(new_n1365), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1331), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n880), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  NOR3_X1   g1171(.A1(new_n1364), .A2(KEYINPUT125), .A3(new_n1310), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1367), .B1(new_n1311), .B2(new_n1366), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1361), .B1(new_n1372), .B2(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1374), .A2(G384), .A3(new_n1331), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1345), .A2(G2897), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1371), .A2(new_n1375), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1376), .B1(new_n1371), .B2(new_n1375), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  AOI22_X1  g1179(.A1(new_n1267), .A2(new_n777), .B1(new_n1280), .B2(new_n1305), .ZN(new_n1380));
  INV_X1    g1180(.A(new_n1277), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1381), .A2(new_n1242), .A3(new_n1312), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1334), .B1(new_n1380), .B2(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1383), .B1(new_n1340), .B2(G378), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1379), .B1(new_n1384), .B2(new_n1345), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT61), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1371), .A2(new_n1375), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1334), .A2(KEYINPUT121), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1215), .A2(new_n1216), .A3(new_n1238), .ZN(new_n1389));
  NAND4_X1  g1189(.A1(new_n1279), .A2(new_n1388), .A3(new_n1389), .A4(new_n1308), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1380), .A2(new_n1382), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(new_n1342), .ZN(new_n1392));
  AOI211_X1 g1192(.A(new_n1345), .B(new_n1387), .C1(new_n1390), .C2(new_n1392), .ZN(new_n1393));
  INV_X1    g1193(.A(KEYINPUT62), .ZN(new_n1394));
  OAI211_X1 g1194(.A(new_n1385), .B(new_n1386), .C1(new_n1393), .C2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1390), .A2(new_n1392), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1396), .A2(new_n1344), .ZN(new_n1397));
  NOR3_X1   g1197(.A1(new_n1397), .A2(KEYINPUT62), .A3(new_n1387), .ZN(new_n1398));
  OAI21_X1  g1198(.A(new_n1360), .B1(new_n1395), .B2(new_n1398), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1400));
  NOR3_X1   g1200(.A1(new_n1349), .A2(KEYINPUT126), .A3(new_n1350), .ZN(new_n1401));
  AOI21_X1  g1201(.A(new_n1355), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1402));
  OAI21_X1  g1202(.A(new_n1400), .B1(new_n1401), .B2(new_n1402), .ZN(new_n1403));
  INV_X1    g1203(.A(KEYINPUT63), .ZN(new_n1404));
  OAI21_X1  g1204(.A(new_n1404), .B1(new_n1397), .B2(new_n1387), .ZN(new_n1405));
  AOI21_X1  g1205(.A(KEYINPUT61), .B1(new_n1397), .B2(new_n1379), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1393), .A2(KEYINPUT63), .ZN(new_n1407));
  NAND4_X1  g1207(.A1(new_n1403), .A2(new_n1405), .A3(new_n1406), .A4(new_n1407), .ZN(new_n1408));
  NAND2_X1  g1208(.A1(new_n1399), .A2(new_n1408), .ZN(G405));
  NAND2_X1  g1209(.A1(G375), .A2(new_n1342), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1410), .A2(new_n1390), .ZN(new_n1411));
  NAND3_X1  g1211(.A1(new_n1411), .A2(new_n1371), .A3(new_n1375), .ZN(new_n1412));
  NAND3_X1  g1212(.A1(new_n1410), .A2(new_n1387), .A3(new_n1390), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1412), .A2(new_n1413), .ZN(new_n1414));
  XNOR2_X1  g1214(.A(new_n1360), .B(new_n1414), .ZN(G402));
endmodule


