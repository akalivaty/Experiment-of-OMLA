//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(G234), .A2(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G952), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G902), .A3(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT21), .B(G898), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(new_n197), .B2(G116), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G116), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(KEYINPUT5), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT84), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(G113), .B1(new_n203), .B2(KEYINPUT5), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(G119), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n198), .B2(new_n201), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(G107), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n217), .A2(G107), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n220), .A2(G104), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n204), .A2(new_n208), .B1(new_n210), .B2(new_n214), .ZN(new_n232));
  INV_X1    g046(.A(new_n228), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n207), .B1(new_n210), .B2(KEYINPUT5), .ZN(new_n235));
  OAI211_X1 g049(.A(KEYINPUT85), .B(new_n228), .C1(new_n216), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G110), .B(G122), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT8), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G224), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G953), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT7), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n251), .A2(KEYINPUT64), .A3(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT64), .B1(new_n251), .B2(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n248), .B(new_n250), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(G143), .B2(new_n247), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n247), .A2(G143), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n256), .A2(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G125), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n247), .B2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n251), .A2(KEYINPUT64), .A3(G146), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n257), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n251), .A2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n248), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n246), .B1(new_n266), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n266), .A2(new_n280), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT7), .B1(new_n242), .B2(KEYINPUT88), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(KEYINPUT88), .B2(new_n242), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n281), .A2(KEYINPUT87), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT78), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n218), .A2(new_n221), .A3(new_n289), .A4(new_n223), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(G101), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n224), .A2(KEYINPUT4), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n202), .A2(new_n203), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n213), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n215), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n288), .A2(new_n298), .A3(G101), .A4(new_n290), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n235), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n233), .A3(new_n215), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(new_n238), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n240), .A2(new_n282), .A3(new_n286), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n304), .A2(KEYINPUT89), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT89), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n297), .A2(new_n299), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n222), .B1(new_n287), .B2(KEYINPUT78), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n292), .B1(new_n311), .B2(new_n290), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n238), .A2(KEYINPUT6), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  INV_X1    g131(.A(new_n238), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT6), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n238), .B1(new_n300), .B2(new_n302), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n316), .A2(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n283), .B(new_n242), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n309), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n317), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n320), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT6), .A3(new_n303), .ZN(new_n328));
  INV_X1    g142(.A(new_n322), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n326), .A2(KEYINPUT83), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G210), .B1(G237), .B2(G902), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n308), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n308), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n187), .B(new_n196), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n251), .A2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n249), .A2(G143), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G134), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n200), .A2(KEYINPUT14), .A3(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(G116), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(G107), .B(new_n341), .C1(new_n343), .C2(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n340), .B(new_n344), .C1(G107), .C2(new_n343), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n337), .B1(new_n346), .B2(KEYINPUT13), .ZN(new_n348));
  OAI21_X1  g162(.A(G134), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n339), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n342), .B(new_n220), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT9), .B(G234), .ZN(new_n354));
  INV_X1    g168(.A(G217), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n354), .A2(new_n355), .A3(G953), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n353), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n305), .ZN(new_n359));
  INV_X1    g173(.A(G478), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n360), .A2(KEYINPUT15), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n359), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT93), .ZN(new_n364));
  NOR2_X1   g178(.A1(G125), .A2(G140), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n265), .B2(G140), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT72), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT72), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n262), .B2(new_n264), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n369), .B(KEYINPUT16), .C1(new_n371), .C2(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n267), .A2(KEYINPUT16), .A3(G140), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(G146), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n247), .B(new_n374), .C1(new_n368), .C2(new_n372), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n364), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n372), .ZN(new_n379));
  INV_X1    g193(.A(new_n365), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n267), .B2(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n369), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n375), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n247), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n373), .A2(G146), .A3(new_n375), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT93), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n189), .A3(G214), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n251), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G131), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n388), .B(G143), .ZN(new_n391));
  INV_X1    g205(.A(G131), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  MUX2_X1   g208(.A(new_n394), .B(new_n390), .S(KEYINPUT17), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n378), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n217), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n247), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n247), .B2(new_n381), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n405), .A2(new_n392), .A3(KEYINPUT90), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n391), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n396), .A2(new_n398), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n398), .B1(new_n396), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n305), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT95), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n305), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT94), .B(G475), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT91), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n390), .A2(new_n393), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n390), .B2(new_n393), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT19), .B1(new_n400), .B2(new_n401), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n381), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT92), .B1(new_n424), .B2(new_n247), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT92), .ZN(new_n426));
  NOR4_X1   g240(.A1(new_n421), .A2(new_n423), .A3(new_n426), .A4(G146), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n420), .B(new_n385), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n408), .ZN(new_n429));
  INV_X1    g243(.A(new_n398), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n396), .A2(new_n398), .A3(new_n408), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT20), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n416), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n335), .A2(new_n363), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n197), .A2(G128), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT70), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n197), .A2(G128), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n197), .A2(KEYINPUT70), .A3(G128), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT24), .B(G110), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n197), .B2(G128), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(G110), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n384), .B2(new_n385), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT73), .B(G110), .Z(new_n458));
  OR2_X1    g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n448), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT74), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n403), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n377), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G137), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n457), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n465), .A2(new_n377), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n455), .B1(new_n376), .B2(new_n377), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT76), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n469), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n470), .B1(new_n457), .B2(new_n466), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n355), .B1(G234), .B2(new_n305), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(KEYINPUT77), .A3(new_n482), .ZN(new_n486));
  INV_X1    g300(.A(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n477), .A3(new_n305), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT25), .A4(new_n305), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n486), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n387), .A2(new_n189), .A3(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G128), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n271), .A2(new_n250), .B1(new_n502), .B2(new_n278), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n339), .B2(G137), .ZN(new_n505));
  INV_X1    g319(.A(G137), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT11), .A3(G134), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n339), .A2(G137), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n392), .A4(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n339), .A2(G137), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n506), .A2(G134), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT65), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n509), .A2(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n260), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G131), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n271), .A2(new_n273), .B1(new_n276), .B2(new_n278), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n297), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n515), .A2(new_n260), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT67), .ZN(new_n526));
  INV_X1    g340(.A(new_n297), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n260), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n522), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n500), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n297), .B1(new_n521), .B2(new_n520), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n499), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n529), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n297), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n530), .A4(new_n498), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n530), .A3(new_n498), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT68), .B(new_n499), .C1(new_n531), .C2(new_n533), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n536), .A2(new_n542), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT32), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n540), .A2(new_n530), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT29), .B1(new_n551), .B2(new_n499), .ZN(new_n552));
  INV_X1    g366(.A(new_n533), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n524), .A2(new_n530), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n498), .B(new_n553), .C1(new_n554), .C2(new_n500), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT69), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT69), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n498), .A2(KEYINPUT29), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n526), .A2(new_n529), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n526), .A2(new_n522), .A3(new_n529), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n561), .A2(new_n532), .B1(new_n562), .B2(new_n297), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n553), .B(new_n560), .C1(new_n563), .C2(new_n500), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n305), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n557), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n494), .B1(new_n550), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G469), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n305), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n260), .A2(KEYINPUT10), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n228), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n233), .A2(new_n260), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n294), .A2(new_n299), .A3(new_n521), .ZN(new_n579));
  INV_X1    g393(.A(new_n502), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n254), .B1(new_n580), .B2(new_n271), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n233), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n520), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n576), .A2(new_n577), .ZN(new_n587));
  INV_X1    g401(.A(new_n520), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n584), .A4(new_n579), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  INV_X1    g405(.A(G227), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n503), .A2(new_n228), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n588), .B1(new_n582), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT80), .A3(KEYINPUT12), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n233), .A2(new_n260), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n502), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n228), .B1(new_n602), .B2(new_n254), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n520), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT80), .B1(new_n598), .B2(KEYINPUT12), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n596), .B(new_n589), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n595), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n573), .B1(new_n610), .B2(new_n572), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n607), .A2(new_n608), .ZN(new_n612));
  INV_X1    g426(.A(new_n589), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n594), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT81), .B1(new_n589), .B2(new_n596), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n589), .A2(new_n596), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT81), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n586), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n614), .B(G469), .C1(new_n615), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n571), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n441), .A2(new_n569), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  AOI21_X1  g436(.A(KEYINPUT77), .B1(new_n480), .B2(new_n482), .ZN(new_n623));
  INV_X1    g437(.A(new_n482), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n484), .B(new_n624), .C1(new_n475), .C2(new_n479), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n623), .A2(new_n625), .A3(new_n492), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n546), .A2(new_n305), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n546), .A2(new_n547), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT96), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(new_n626), .A3(new_n634), .A4(new_n620), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n359), .A2(new_n360), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT33), .B1(new_n356), .B2(KEYINPUT97), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n358), .B(new_n640), .Z(new_n641));
  NOR2_X1   g455(.A1(new_n360), .A2(G902), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n638), .A2(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n416), .B2(new_n439), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT99), .B1(new_n645), .B2(new_n335), .ZN(new_n646));
  INV_X1    g460(.A(new_n335), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n644), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n636), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(new_n415), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n411), .B2(KEYINPUT95), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n414), .B1(new_n436), .B2(new_n438), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n363), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n335), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n457), .A2(new_n466), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n482), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n493), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n620), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n631), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n441), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(G472), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n565), .B1(new_n556), .B2(KEYINPUT69), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n672), .B1(new_n673), .B2(new_n559), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n548), .A3(new_n549), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n187), .B1(new_n333), .B2(new_n334), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n667), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT100), .B(G900), .Z(new_n679));
  AOI21_X1  g493(.A(new_n191), .B1(new_n679), .B2(new_n193), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n362), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n416), .A2(new_n439), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n678), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT102), .B(G128), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G30));
  NOR2_X1   g502(.A1(new_n333), .A2(new_n334), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n363), .A2(new_n187), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n690), .A2(new_n655), .A3(new_n666), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n680), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n620), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n694), .A2(new_n695), .ZN(new_n698));
  OR3_X1    g512(.A1(new_n697), .A2(KEYINPUT40), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT40), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT32), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n630), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n562), .A2(new_n297), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n530), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n499), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n543), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n305), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n702), .A2(new_n703), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT104), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n702), .A2(new_n714), .A3(new_n711), .A4(new_n703), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n692), .A2(new_n699), .A3(new_n700), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  INV_X1    g533(.A(new_n680), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n644), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n719), .B1(new_n721), .B2(new_n676), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n675), .A2(new_n667), .ZN(new_n723));
  INV_X1    g537(.A(new_n187), .ZN(new_n724));
  INV_X1    g538(.A(new_n332), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n323), .A2(new_n330), .ZN(new_n726));
  INV_X1    g540(.A(new_n307), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n304), .A2(KEYINPUT89), .A3(new_n305), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n308), .A2(new_n331), .A3(new_n332), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n724), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n644), .A2(new_n732), .A3(KEYINPUT106), .A4(new_n720), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n722), .A2(new_n723), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NAND2_X1  g549(.A1(new_n702), .A2(new_n703), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n626), .B1(new_n736), .B2(new_n674), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n610), .A2(new_n572), .ZN(new_n738));
  INV_X1    g552(.A(new_n609), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n596), .B1(new_n586), .B2(new_n589), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n572), .B(new_n305), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n738), .A2(new_n742), .A3(new_n571), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n646), .A2(new_n745), .A3(new_n649), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n657), .A2(new_n569), .A3(new_n743), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  AND3_X1   g564(.A1(new_n743), .A2(new_n196), .A3(new_n666), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n677), .A2(new_n362), .A3(new_n655), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  OAI21_X1  g567(.A(new_n553), .B1(new_n563), .B2(new_n500), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n499), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n544), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n542), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n755), .B2(new_n544), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n547), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT108), .B(G472), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n628), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n626), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n689), .A2(new_n655), .A3(new_n691), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n744), .A2(new_n195), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NAND2_X1  g581(.A1(new_n730), .A2(new_n731), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n187), .A3(new_n743), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n655), .A2(new_n643), .A3(new_n680), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n666), .A2(new_n760), .A3(new_n762), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT109), .B(G125), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G27));
  INV_X1    g589(.A(new_n573), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n619), .A2(new_n741), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n570), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n780), .A3(new_n570), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n689), .A3(new_n187), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n720), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n703), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n546), .A2(KEYINPUT111), .A3(KEYINPUT32), .A4(new_n547), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n568), .A2(new_n786), .A3(new_n702), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n626), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n788), .B2(new_n626), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n784), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n730), .A2(new_n187), .A3(new_n731), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n780), .B1(new_n777), .B2(new_n570), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n569), .A2(new_n797), .A3(new_n781), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n794), .B1(new_n798), .B2(new_n721), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n684), .A2(new_n685), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n684), .A2(new_n685), .ZN(new_n805));
  INV_X1    g619(.A(new_n782), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(KEYINPUT113), .A4(new_n569), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  OAI21_X1  g623(.A(new_n614), .B1(new_n615), .B2(new_n618), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n572), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n573), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n741), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n570), .B(new_n693), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n795), .B(KEYINPUT114), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n631), .A2(new_n666), .ZN(new_n820));
  INV_X1    g634(.A(new_n643), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n655), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT43), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n655), .A2(KEYINPUT43), .A3(new_n821), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n818), .B(new_n819), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  OAI21_X1  g645(.A(new_n570), .B1(new_n815), .B2(new_n816), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(KEYINPUT47), .B(new_n570), .C1(new_n815), .C2(new_n816), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n675), .A2(new_n187), .A3(new_n689), .A4(new_n494), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n837), .A2(new_n838), .A3(new_n721), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n837), .B2(new_n721), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n666), .A2(new_n778), .A3(new_n680), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n716), .A2(new_n764), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n686), .A2(new_n845), .A3(new_n773), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n733), .A2(new_n723), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT106), .B1(new_n771), .B2(new_n732), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n843), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(KEYINPUT117), .B(new_n843), .C1(new_n846), .C2(new_n849), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n772), .A2(new_n644), .A3(new_n720), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n675), .A2(new_n667), .A3(new_n676), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n770), .A2(new_n854), .B1(new_n805), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n845), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n416), .A2(new_n439), .A3(new_n362), .A4(new_n720), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n795), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n620), .B(new_n666), .C1(new_n736), .C2(new_n674), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n860), .B2(KEYINPUT116), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n861), .A2(new_n863), .B1(new_n854), .B2(new_n806), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n800), .A2(new_n808), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n749), .A2(new_n766), .A3(new_n669), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n621), .A2(new_n752), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n645), .A2(new_n656), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n632), .A2(new_n868), .A3(new_n647), .A4(new_n635), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n746), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n858), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n800), .A2(new_n808), .A3(new_n864), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n857), .A2(new_n850), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n869), .A2(new_n621), .A3(new_n752), .ZN(new_n875));
  INV_X1    g689(.A(new_n746), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n749), .A2(new_n766), .A3(new_n669), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(KEYINPUT53), .A2(new_n873), .A3(new_n874), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n799), .A2(new_n793), .B1(new_n804), .B2(new_n807), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n882), .A3(new_n864), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n857), .A2(new_n850), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n858), .A2(KEYINPUT53), .A3(new_n871), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n744), .A2(new_n795), .A3(new_n494), .A4(new_n190), .ZN(new_n889));
  INV_X1    g703(.A(new_n716), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n655), .A4(new_n643), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n190), .B1(new_n824), .B2(new_n825), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n744), .A2(new_n795), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n772), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n690), .A2(new_n724), .A3(new_n743), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n892), .A3(KEYINPUT50), .A4(new_n763), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT50), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n763), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n819), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT118), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n892), .A2(new_n819), .A3(new_n906), .A4(new_n763), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n738), .A2(new_n742), .A3(new_n570), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n905), .B(new_n907), .C1(new_n836), .C2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n903), .A2(new_n909), .A3(KEYINPUT51), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT51), .B1(new_n903), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n892), .A2(new_n763), .A3(new_n770), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n889), .A2(new_n890), .A3(new_n644), .ZN(new_n913));
  AND4_X1   g727(.A1(G952), .A2(new_n912), .A3(new_n189), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n894), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT48), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n789), .B(KEYINPUT112), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n910), .A2(new_n911), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n880), .A2(new_n888), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(G952), .A2(G953), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT119), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n738), .A2(new_n742), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT49), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n626), .A2(new_n187), .A3(new_n570), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n822), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n890), .A3(new_n690), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G75));
  AOI21_X1  g749(.A(new_n305), .B1(new_n885), .B2(new_n886), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(G210), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n321), .B(new_n322), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n189), .A2(G952), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G51));
  NAND2_X1  g759(.A1(new_n885), .A2(new_n886), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n888), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n573), .B(KEYINPUT57), .Z(new_n950));
  OAI22_X1  g764(.A1(new_n949), .A2(new_n950), .B1(new_n740), .B2(new_n739), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n812), .A2(new_n813), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT121), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n936), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n944), .B1(new_n951), .B2(new_n954), .ZN(G54));
  AND2_X1   g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n936), .A2(new_n433), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n433), .B1(new_n936), .B2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n944), .ZN(G60));
  NAND2_X1  g773(.A1(new_n880), .A2(new_n888), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT59), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n641), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n641), .A2(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n944), .B1(new_n948), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n944), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n641), .B1(new_n960), .B2(new_n962), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT122), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n969), .A2(new_n976), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT60), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n946), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n479), .A3(new_n475), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n946), .A2(new_n664), .A3(new_n979), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n973), .A4(new_n982), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G66));
  OAI21_X1  g801(.A(G953), .B1(new_n194), .B2(new_n241), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n878), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n321), .B1(G898), .B2(new_n189), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  NAND3_X1  g805(.A1(new_n917), .A2(new_n818), .A3(new_n764), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n856), .A2(new_n734), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n882), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n993), .A2(new_n995), .A3(new_n830), .A4(new_n841), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n538), .A2(new_n539), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT123), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n424), .ZN(new_n1000));
  INV_X1    g814(.A(G900), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n189), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1004));
  NOR2_X1   g818(.A1(new_n737), .A2(new_n795), .ZN(new_n1005));
  INV_X1    g819(.A(new_n698), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n696), .A4(new_n868), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n830), .A2(new_n841), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n994), .A2(new_n717), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n994), .A2(new_n717), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1004), .B1(new_n1013), .B2(new_n189), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1003), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(G953), .B1(new_n592), .B2(new_n1001), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n996), .B2(new_n870), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n551), .A2(new_n498), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n944), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n551), .A2(new_n498), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1019), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1024), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n872), .B2(new_n879), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1008), .A2(new_n1010), .A3(new_n878), .A4(new_n1012), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1031), .A2(new_n1019), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1030), .B1(new_n1032), .B2(new_n1023), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1031), .A2(new_n1019), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1034), .A2(KEYINPUT126), .A3(new_n1024), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1028), .A2(new_n1029), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1033), .A2(new_n1027), .A3(new_n1022), .A4(new_n1035), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT127), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n1038), .ZN(G57));
endmodule


