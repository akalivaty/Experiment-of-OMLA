//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g0011(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G97), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n205), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n208), .B(new_n219), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(G97), .B(G107), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n221), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n246), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G283), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G97), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n215), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n211), .A2(new_n212), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G116), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n259), .A4(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n264), .A2(new_n265), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(G1), .B2(new_n255), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G116), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT78), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(KEYINPUT78), .A3(G116), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT5), .B(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n255), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n278), .A2(new_n280), .A3(G274), .A4(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n282), .B2(new_n278), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(G270), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G303), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n289), .B(new_n294), .C1(new_n296), .C2(new_n230), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n213), .B1(new_n255), .B2(new_n279), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n277), .B1(G200), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n287), .A2(G190), .A3(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n287), .B2(new_n300), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(KEYINPUT21), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n287), .A2(G179), .A3(new_n300), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n277), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT21), .B1(new_n277), .B2(new_n306), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(KEYINPUT79), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT79), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n313), .B(KEYINPUT21), .C1(new_n277), .C2(new_n306), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n304), .B(new_n310), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G58), .A2(G68), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT67), .B(G58), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(G68), .ZN(new_n319));
  INV_X1    g0119(.A(G20), .ZN(new_n320));
  INV_X1    g0120(.A(G159), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G20), .A2(G33), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n319), .A2(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n290), .A2(G33), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n320), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n221), .B1(new_n328), .B2(KEYINPUT7), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n293), .A2(new_n215), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT71), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT7), .B1(new_n288), .B2(G20), .ZN(new_n333));
  AND4_X1   g0133(.A1(KEYINPUT71), .A2(new_n333), .A3(new_n331), .A4(G68), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n325), .C1(new_n332), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n320), .A2(KEYINPUT65), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT65), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n330), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n290), .A3(G33), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n292), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n328), .A2(new_n330), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n221), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n336), .B1(new_n348), .B2(new_n324), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n335), .A2(new_n259), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT8), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G58), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n318), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n268), .ZN(new_n354));
  INV_X1    g0154(.A(new_n259), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G1), .B2(new_n320), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n356), .B2(new_n353), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n350), .A2(KEYINPUT73), .A3(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n363));
  INV_X1    g0163(.A(G274), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n280), .A2(new_n363), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n228), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G223), .A2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G226), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n288), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n255), .B2(new_n223), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n373), .B2(new_n299), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G179), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n305), .B2(new_n374), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n361), .A2(new_n362), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT18), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  AOI21_X1  g0180(.A(G20), .B1(new_n291), .B2(new_n292), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n381), .B2(new_n330), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n337), .A2(new_n339), .A3(new_n330), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n288), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n333), .A2(new_n331), .A3(KEYINPUT71), .A4(G68), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n324), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n355), .B1(new_n387), .B2(KEYINPUT16), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n357), .B1(new_n388), .B2(new_n349), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n374), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G200), .B2(new_n374), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n379), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n379), .A2(new_n350), .A3(new_n358), .A4(new_n392), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT17), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n350), .A2(new_n392), .A3(new_n358), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n361), .A2(new_n399), .A3(new_n362), .A4(new_n376), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n378), .A2(new_n395), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n268), .A2(new_n247), .ZN(new_n402));
  INV_X1    g0202(.A(G150), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n323), .B1(new_n201), .B2(new_n320), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n215), .A2(G33), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n406), .B2(new_n353), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n402), .B1(new_n356), .B2(new_n247), .C1(new_n407), .C2(new_n355), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT9), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n366), .B1(new_n367), .B2(new_n370), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n288), .A2(G222), .A3(new_n295), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n288), .A2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(G223), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n411), .B1(new_n202), .B2(new_n288), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n414), .B2(new_n299), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G190), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(KEYINPUT10), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(KEYINPUT10), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n408), .B1(new_n415), .B2(G169), .ZN(new_n423));
  INV_X1    g0223(.A(G179), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n415), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(new_n296), .C2(new_n370), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n299), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n280), .A2(new_n363), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT68), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT68), .ZN(new_n435));
  OAI21_X1  g0235(.A(G238), .B1(new_n367), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n366), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n434), .A2(new_n436), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n431), .A4(new_n366), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n441), .A3(G190), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT69), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n268), .A2(new_n221), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n221), .B2(new_n356), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT11), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n322), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n405), .B2(new_n202), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n259), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n448), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n438), .A2(new_n441), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(G200), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n438), .B2(new_n441), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT14), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(new_n454), .B2(new_n424), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n459), .A2(new_n460), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT15), .B(G87), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n406), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n227), .A2(KEYINPUT8), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n352), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n322), .B1(new_n340), .B2(G77), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n355), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n268), .A2(new_n202), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n356), .B2(new_n202), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G107), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n412), .A2(new_n222), .B1(new_n475), .B2(new_n288), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n293), .A2(new_n228), .A3(G1698), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n299), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n365), .B1(new_n433), .B2(G244), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n474), .B1(new_n480), .B2(G200), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n390), .B2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n305), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n424), .A3(new_n479), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n401), .A2(new_n427), .A3(new_n464), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  INV_X1    g0288(.A(G244), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n296), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n295), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n490), .A2(new_n254), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n299), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n286), .A2(G257), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n283), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n305), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n475), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n245), .B2(KEYINPUT6), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n340), .B1(G77), .B2(new_n322), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n341), .A2(new_n345), .B1(new_n328), .B2(new_n330), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n475), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n259), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n267), .A2(G97), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n271), .B2(G97), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n496), .B1(new_n493), .B2(new_n299), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n424), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n499), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n507), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n504), .B2(new_n259), .ZN(new_n513));
  AOI211_X1 g0313(.A(G190), .B(new_n496), .C1(new_n299), .C2(new_n493), .ZN(new_n514));
  AOI21_X1  g0314(.A(G200), .B1(new_n494), .B2(new_n497), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n215), .A2(new_n288), .A3(G87), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT23), .A2(G107), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G20), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT23), .A2(G107), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n340), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n520), .B1(new_n519), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n259), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n288), .A2(G250), .A3(new_n295), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(new_n412), .C2(new_n230), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n299), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n286), .A2(G264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n283), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n416), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n531), .A2(new_n299), .B1(new_n286), .B2(G264), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n390), .A3(new_n283), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT25), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n267), .B2(G107), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n475), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n271), .A2(G107), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n528), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n528), .A2(new_n538), .A3(KEYINPUT80), .A4(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n517), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n405), .B2(new_n229), .ZN(new_n549));
  OR2_X1    g0349(.A1(KEYINPUT75), .A2(G87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT75), .A2(G87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n229), .A3(new_n475), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n429), .A2(new_n548), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n340), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n215), .A2(new_n288), .A3(G68), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n549), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n355), .B1(new_n556), .B2(KEYINPUT76), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT76), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n549), .A2(new_n554), .A3(new_n558), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n465), .A2(new_n268), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n271), .A2(new_n466), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT77), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n280), .B(G250), .C1(G1), .C2(new_n281), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n282), .A2(G274), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n288), .A2(G244), .A3(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n296), .C2(new_n222), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n299), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n305), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n424), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n564), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n557), .A2(new_n559), .B1(new_n268), .B2(new_n465), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(G200), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n271), .A2(G87), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n534), .A2(new_n305), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G179), .B2(new_n534), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n528), .B2(new_n542), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n316), .A2(new_n487), .A3(new_n547), .A4(new_n585), .ZN(G372));
  NAND2_X1  g0386(.A1(new_n528), .A2(new_n542), .ZN(new_n587));
  INV_X1    g0387(.A(new_n583), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n310), .C1(new_n312), .C2(new_n314), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n570), .A2(new_n591), .A3(new_n299), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n570), .B2(new_n299), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n566), .B(new_n565), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(new_n576), .A3(new_n577), .A4(new_n579), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n305), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n564), .A2(new_n597), .A3(new_n574), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n547), .A2(new_n590), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT26), .B1(new_n581), .B2(new_n511), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  INV_X1    g0403(.A(new_n511), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n598), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n487), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n395), .A2(new_n398), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n485), .A2(KEYINPUT82), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n483), .A2(new_n474), .A3(new_n610), .A4(new_n484), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n456), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n608), .B1(new_n612), .B2(new_n463), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n359), .A2(new_n376), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n614), .B(KEYINPUT18), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n422), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n607), .A2(new_n426), .A3(new_n616), .ZN(G369));
  NAND2_X1  g0417(.A1(new_n316), .A2(KEYINPUT83), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n215), .A2(new_n266), .A3(G13), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  OAI21_X1  g0420(.A(G213), .B1(new_n619), .B2(KEYINPUT27), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n277), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n315), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n310), .B1(new_n312), .B2(new_n314), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n618), .A2(new_n627), .B1(new_n628), .B2(new_n625), .ZN(new_n629));
  INV_X1    g0429(.A(G330), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n624), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n584), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n545), .A2(new_n546), .B1(new_n587), .B2(new_n624), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n584), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n636), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n628), .A2(new_n633), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(G399));
  INV_X1    g0443(.A(KEYINPUT84), .ZN(new_n644));
  INV_X1    g0444(.A(new_n206), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(G41), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n206), .A2(KEYINPUT84), .A3(new_n279), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n552), .A2(G116), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G1), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n217), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT28), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n599), .B2(new_n511), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n604), .A2(new_n603), .A3(new_n575), .A4(new_n580), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n601), .A2(new_n598), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n633), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT29), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n606), .A2(new_n633), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(KEYINPUT29), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n316), .A2(new_n547), .A3(new_n585), .A4(new_n633), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT31), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT85), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n494), .A2(new_n536), .A3(new_n497), .A4(new_n571), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n308), .ZN(new_n665));
  AOI21_X1  g0465(.A(G179), .B1(new_n287), .B2(new_n300), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n594), .A2(new_n534), .A3(new_n498), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n663), .B1(new_n664), .B2(new_n308), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n536), .A2(new_n571), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n309), .A2(new_n670), .A3(KEYINPUT30), .A4(new_n509), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n662), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n661), .B1(new_n673), .B2(new_n633), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n660), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n659), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n652), .B1(new_n680), .B2(G1), .ZN(G364));
  AND2_X1   g0481(.A1(new_n215), .A2(G13), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G45), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT86), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n266), .B1(new_n683), .B2(KEYINPUT86), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n648), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n631), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n629), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(G330), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n645), .A2(new_n293), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(G355), .B1(new_n260), .B2(new_n645), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n252), .A2(new_n281), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n645), .A2(new_n288), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(G45), .B2(new_n217), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n214), .B1(G20), .B2(new_n305), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G13), .A2(G33), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G20), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n697), .B2(KEYINPUT87), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n688), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  NOR4_X1   g0505(.A1(new_n215), .A2(G179), .A3(G190), .A4(new_n416), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n215), .A2(new_n424), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n390), .A2(new_n416), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT92), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(G283), .A2(new_n710), .B1(new_n715), .B2(G326), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n390), .A2(G179), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n215), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G294), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n293), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR4_X1   g0520(.A1(new_n215), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(G329), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n712), .A2(G20), .A3(new_n424), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT90), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n390), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n711), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n728), .A2(G303), .B1(new_n731), .B2(G322), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n711), .A2(new_n390), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n416), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  AOI22_X1  g0536(.A1(G311), .A2(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n716), .A2(new_n722), .A3(new_n732), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n318), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n288), .B1(new_n229), .B2(new_n718), .C1(new_n730), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n550), .A2(new_n551), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n727), .A2(new_n742), .B1(new_n713), .B2(new_n247), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n740), .B(new_n743), .C1(G68), .C2(new_n735), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n721), .A2(G159), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT89), .B(KEYINPUT32), .Z(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n710), .A2(G107), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n734), .A2(KEYINPUT88), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n734), .A2(KEYINPUT88), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n202), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n738), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  AOI21_X1  g0555(.A(new_n705), .B1(new_n755), .B2(new_n699), .ZN(new_n756));
  INV_X1    g0556(.A(new_n702), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n690), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n691), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(G396));
  NAND2_X1  g0560(.A1(new_n474), .A2(new_n624), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n482), .A2(new_n485), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n609), .A2(new_n474), .A3(new_n611), .A4(new_n624), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n658), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n764), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n606), .A2(new_n633), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n688), .B1(new_n768), .B2(new_n678), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n678), .B2(new_n768), .ZN(new_n770));
  INV_X1    g0570(.A(new_n699), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n701), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n688), .B1(G77), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  INV_X1    g0574(.A(new_n752), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G116), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n710), .A2(G87), .ZN(new_n777));
  INV_X1    g0577(.A(new_n721), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(new_n719), .B2(new_n730), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G107), .B2(new_n728), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n293), .B1(new_n229), .B2(new_n718), .C1(new_n713), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G283), .B2(new_n735), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n727), .A2(new_n247), .ZN(new_n786));
  INV_X1    g0586(.A(G132), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n288), .B1(new_n739), .B2(new_n718), .C1(new_n778), .C2(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n710), .C2(G68), .ZN(new_n789));
  INV_X1    g0589(.A(new_n713), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G137), .A2(new_n790), .B1(new_n731), .B2(G143), .ZN(new_n791));
  INV_X1    g0591(.A(new_n735), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n403), .B2(new_n792), .C1(new_n752), .C2(new_n321), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n789), .B1(new_n794), .B2(KEYINPUT34), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT34), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n785), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n774), .B1(new_n798), .B2(new_n699), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n766), .B2(new_n701), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n770), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G384));
  OR2_X1    g0602(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n803), .A2(G116), .A3(new_n216), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT36), .Z(new_n806));
  OAI211_X1 g0606(.A(G77), .B(new_n218), .C1(new_n739), .C2(new_n221), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n266), .B(G13), .C1(new_n807), .C2(new_n248), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n615), .A2(new_n622), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n485), .A2(new_n624), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n767), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n453), .A2(new_n624), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n456), .A2(new_n463), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n453), .B(new_n624), .C1(new_n461), .C2(new_n462), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n388), .B1(KEYINPUT16), .B2(new_n387), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n622), .B1(new_n818), .B2(new_n358), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n401), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n389), .A2(new_n379), .A3(new_n392), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n622), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n376), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n358), .B2(new_n818), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n376), .A2(new_n824), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n361), .A2(new_n362), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n821), .A2(new_n822), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n820), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT38), .B1(new_n820), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n810), .B1(new_n817), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT95), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n820), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT96), .B1(new_n830), .B2(new_n832), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n361), .A2(new_n362), .A3(new_n824), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n614), .A2(new_n396), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n393), .A2(new_n394), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT96), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(new_n831), .A4(new_n829), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n841), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n842), .B1(new_n608), .B2(new_n615), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n850), .B2(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n463), .A2(new_n624), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT95), .B(new_n810), .C1(new_n817), .C2(new_n836), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n839), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n616), .A2(new_n426), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n659), .B2(new_n487), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n859), .B(new_n861), .Z(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n672), .A2(new_n669), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT31), .B(new_n624), .C1(new_n864), .C2(new_n668), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n660), .A2(new_n674), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n764), .B1(new_n814), .B2(new_n815), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n834), .B2(new_n835), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n866), .A2(KEYINPUT40), .A3(new_n867), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n863), .A2(new_n869), .B1(new_n851), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n487), .A3(new_n866), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n487), .B2(new_n866), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n862), .A2(new_n875), .B1(new_n266), .B2(new_n682), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n862), .A2(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n809), .B1(new_n879), .B2(new_n880), .ZN(G367));
  INV_X1    g0681(.A(new_n238), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n695), .ZN(new_n883));
  INV_X1    g0683(.A(new_n703), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n645), .B2(new_n466), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n687), .B(new_n686), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT104), .Z(new_n887));
  AOI21_X1  g0687(.A(new_n633), .B1(new_n576), .B2(new_n579), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n574), .A3(new_n564), .A4(new_n597), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n599), .B2(new_n888), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n728), .A2(KEYINPUT46), .A3(G116), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT46), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n727), .B2(new_n260), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n891), .B(new_n893), .C1(new_n719), .C2(new_n792), .ZN(new_n894));
  INV_X1    g0694(.A(G317), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n293), .B1(new_n475), .B2(new_n718), .C1(new_n778), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(G303), .B2(new_n731), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n710), .A2(G97), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT105), .B(G311), .Z(new_n899));
  OAI211_X1 g0699(.A(new_n897), .B(new_n898), .C1(new_n714), .C2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n894), .B(new_n900), .C1(G283), .C2(new_n775), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT106), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n730), .A2(new_n403), .B1(new_n221), .B2(new_n718), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n715), .A2(G143), .B1(KEYINPUT107), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n710), .A2(G77), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(new_n905), .C1(KEYINPUT107), .C2(new_n903), .ZN(new_n906));
  INV_X1    g0706(.A(G137), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n288), .B1(new_n778), .B2(new_n907), .C1(new_n727), .C2(new_n739), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G159), .B2(new_n735), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n247), .B2(new_n752), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n913));
  AND2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n699), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n887), .B1(new_n757), .B2(new_n890), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n604), .A2(new_n624), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n511), .B(new_n516), .C1(new_n513), .C2(new_n633), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n642), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT45), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n642), .A2(new_n919), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(KEYINPUT101), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(KEYINPUT101), .ZN(new_n925));
  XNOR2_X1  g0725(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n921), .B(new_n927), .C1(new_n924), .C2(new_n926), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(new_n637), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n637), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n631), .A2(KEYINPUT103), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT102), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n639), .B2(new_n640), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n641), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n680), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n680), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n648), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n686), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n890), .A2(KEYINPUT98), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n890), .A2(KEYINPUT98), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n936), .A2(new_n919), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT99), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(KEYINPUT99), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(KEYINPUT42), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n511), .B1(new_n918), .B2(new_n589), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n633), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT42), .B1(new_n949), .B2(new_n950), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n946), .B(new_n956), .C1(KEYINPUT43), .C2(new_n890), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n946), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n637), .A2(new_n919), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n916), .B1(new_n943), .B2(new_n960), .ZN(G387));
  OAI21_X1  g0761(.A(new_n695), .B1(new_n242), .B2(new_n281), .ZN(new_n962));
  INV_X1    g0762(.A(new_n692), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n649), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n469), .A2(new_n247), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n966));
  AOI21_X1  g0766(.A(G45), .B1(G68), .B2(G77), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n966), .A2(new_n649), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n964), .A2(new_n969), .B1(new_n475), .B2(new_n645), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n728), .A2(G77), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n288), .C1(new_n465), .C2(new_n718), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n353), .B2(new_n735), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n734), .A2(G68), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n247), .A2(new_n730), .B1(new_n713), .B2(new_n321), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G150), .B2(new_n721), .ZN(new_n976));
  AND4_X1   g0776(.A1(new_n898), .A2(new_n973), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G322), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n714), .A2(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n792), .A2(new_n899), .B1(new_n730), .B2(new_n895), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n775), .C2(G303), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT48), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT48), .ZN(new_n983));
  INV_X1    g0783(.A(new_n718), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n728), .A2(G294), .B1(G283), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT49), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n288), .B1(new_n721), .B2(G326), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n260), .B2(new_n709), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n987), .B2(KEYINPUT49), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n977), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n688), .B1(new_n884), .B2(new_n970), .C1(new_n992), .C2(new_n771), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n636), .B2(new_n702), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n937), .B2(new_n686), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n938), .A2(new_n687), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n937), .A2(new_n680), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G393));
  NAND2_X1  g0798(.A1(new_n775), .A2(new_n469), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n293), .B1(new_n984), .B2(G77), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n721), .A2(G143), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n727), .C2(new_n221), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G50), .B2(new_n735), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n403), .A2(new_n713), .B1(new_n730), .B2(new_n321), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT51), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n999), .A2(new_n1003), .A3(new_n777), .A4(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n293), .B1(new_n260), .B2(new_n718), .C1(new_n778), .C2(new_n978), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G283), .B2(new_n728), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n779), .A2(new_n730), .B1(new_n713), .B2(new_n895), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT52), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G294), .A2(new_n734), .B1(new_n735), .B2(G303), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n748), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n771), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n246), .A2(new_n695), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n703), .C1(new_n229), .C2(new_n206), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT109), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n688), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n919), .B2(new_n757), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n686), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n931), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n931), .A2(new_n938), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n939), .A2(new_n687), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT110), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT110), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n939), .A2(new_n1027), .A3(new_n687), .A4(new_n1024), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1023), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G390));
  NAND3_X1  g0830(.A1(new_n655), .A2(new_n633), .A3(new_n766), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n811), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n856), .B1(new_n1032), .B2(new_n816), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n851), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n679), .A2(new_n867), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n853), .A2(new_n854), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n856), .B1(new_n812), .B2(new_n816), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1034), .B(new_n1035), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n866), .A2(G330), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n867), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n853), .B2(new_n854), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1033), .A2(new_n851), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n816), .B1(new_n679), .B2(new_n766), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n812), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n816), .B1(new_n1039), .B2(new_n766), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1035), .A2(new_n811), .A3(new_n1031), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1039), .A2(new_n487), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n861), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n648), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1038), .A2(new_n1044), .A3(new_n1052), .A4(new_n1050), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n688), .B1(new_n353), .B2(new_n772), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT54), .B(G143), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n775), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n721), .A2(G125), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n787), .B2(new_n730), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n288), .B1(new_n321), .B2(new_n718), .C1(new_n713), .C2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(G137), .C2(new_n735), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n727), .A2(new_n403), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n710), .A2(G50), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1060), .A2(new_n1065), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n752), .A2(new_n229), .B1(new_n475), .B2(new_n792), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT111), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n730), .A2(new_n260), .B1(new_n202), .B2(new_n718), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT112), .Z(new_n1073));
  INV_X1    g0873(.A(G283), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n293), .B1(new_n713), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n727), .A2(new_n223), .B1(new_n778), .B2(new_n719), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n710), .C2(G68), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1071), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1070), .A2(KEYINPUT111), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1069), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1057), .B1(new_n1080), .B2(new_n699), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1036), .B2(new_n701), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1056), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G378));
  NAND2_X1  g0885(.A1(new_n1055), .A2(new_n1052), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT38), .B1(new_n848), .B2(new_n849), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n870), .B1(new_n834), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n866), .A2(new_n867), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n820), .A2(new_n833), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT38), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1092), .B2(new_n840), .ZN(new_n1093));
  OAI211_X1 g0893(.A(G330), .B(new_n1088), .C1(new_n1093), .C2(KEYINPUT40), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n408), .A2(new_n824), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n427), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n427), .A2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1099), .A3(new_n1095), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1094), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT114), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1094), .A2(KEYINPUT114), .A3(new_n1106), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n859), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n869), .A2(new_n863), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1113), .A2(G330), .A3(new_n1088), .A4(new_n1105), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n871), .A2(KEYINPUT115), .A3(G330), .A4(new_n1105), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1111), .A2(new_n1112), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1112), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1120));
  OAI211_X1 g0920(.A(KEYINPUT57), .B(new_n1086), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1086), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1094), .A2(KEYINPUT114), .A3(new_n1106), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT114), .B1(new_n1094), .B2(new_n1106), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1127), .A2(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n859), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1111), .A2(new_n1112), .A3(new_n1118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n1086), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1123), .A2(new_n1126), .A3(new_n1135), .A4(new_n687), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1106), .A2(new_n700), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n688), .B1(G50), .B2(new_n772), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT113), .Z(new_n1139));
  AOI211_X1 g0939(.A(G41), .B(new_n288), .C1(new_n984), .C2(G68), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n971), .B(new_n1140), .C1(new_n229), .C2(new_n792), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n709), .A2(new_n739), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G107), .A2(new_n731), .B1(new_n790), .B2(G116), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n1074), .C2(new_n778), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1141), .B(new_n1145), .C1(new_n466), .C2(new_n734), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1146), .A2(KEYINPUT58), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n731), .A2(G128), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n790), .A2(G125), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n403), .B2(new_n718), .C1(new_n727), .C2(new_n1058), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n734), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n787), .A2(new_n792), .B1(new_n1152), .B2(new_n907), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n710), .A2(G159), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n721), .C2(G124), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1146), .A2(KEYINPUT58), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n279), .B1(new_n290), .B2(new_n255), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n247), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1147), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1139), .B1(new_n1164), .B2(new_n699), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1134), .A2(new_n686), .B1(new_n1137), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1136), .A2(new_n1166), .ZN(G375));
  OAI21_X1  g0967(.A(new_n688), .B1(G68), .B2(new_n772), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n816), .A2(new_n701), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n288), .B1(new_n247), .B2(new_n718), .C1(new_n727), .C2(new_n321), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G150), .B2(new_n734), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n735), .A2(new_n1059), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n787), .A2(new_n713), .B1(new_n730), .B2(new_n907), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G128), .B2(new_n721), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1143), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n752), .A2(new_n475), .B1(new_n260), .B2(new_n792), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT117), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n293), .B1(new_n718), .B2(new_n465), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G303), .B2(new_n721), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n727), .A2(new_n229), .B1(new_n730), .B2(new_n1074), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G294), .B2(new_n790), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n905), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1176), .A2(KEYINPUT117), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1175), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1168), .B(new_n1169), .C1(new_n699), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1050), .B2(new_n686), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT118), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n942), .A3(new_n1053), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(G381));
  INV_X1    g0990(.A(G387), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(G375), .A2(G378), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n1029), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT119), .ZN(G407));
  INV_X1    g0995(.A(new_n1192), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n623), .A2(G213), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT120), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G407), .B(G213), .C1(new_n1196), .C2(new_n1198), .ZN(G409));
  INV_X1    g0999(.A(KEYINPUT127), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1136), .A2(G378), .A3(new_n1166), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1136), .A2(G378), .A3(KEYINPUT121), .A4(new_n1166), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT122), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1124), .B2(new_n941), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1134), .A2(KEYINPUT122), .A3(new_n942), .A4(new_n1086), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1166), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1084), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1205), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1198), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1188), .A2(KEYINPUT124), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT60), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1053), .A2(new_n687), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1187), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(new_n801), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n801), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT62), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1212), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1211), .A2(KEYINPUT123), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1210), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT123), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1223), .A2(new_n1198), .A3(new_n1227), .A4(new_n1220), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G2897), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1198), .A2(new_n1231), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1219), .B(new_n1232), .Z(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT61), .B1(new_n1212), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1200), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1212), .A2(new_n1221), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1198), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1238));
  AOI211_X1 g1038(.A(KEYINPUT123), .B(new_n1224), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1219), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1237), .B1(new_n1240), .B2(KEYINPUT62), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(KEYINPUT127), .A3(new_n1234), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G387), .A2(new_n1029), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1029), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(new_n759), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(KEYINPUT126), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1245), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT126), .B1(G387), .B2(new_n1029), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1246), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1248), .A2(new_n1243), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1236), .A2(new_n1242), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1211), .A2(KEYINPUT63), .A3(new_n1198), .A4(new_n1220), .ZN(new_n1255));
  AND4_X1   g1055(.A1(new_n1254), .A2(new_n1247), .A3(new_n1251), .A4(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1223), .A2(new_n1198), .A3(new_n1227), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1233), .A3(KEYINPUT125), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1233), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1256), .B1(KEYINPUT63), .B2(new_n1240), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1253), .A2(new_n1261), .ZN(G405));
  AOI22_X1  g1062(.A1(new_n1203), .A2(new_n1204), .B1(new_n1084), .B2(G375), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n1219), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1252), .B(new_n1264), .ZN(G402));
endmodule


