//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G134), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G137), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n187), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n198), .B1(new_n203), .B2(G143), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n205), .B1(new_n203), .B2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n196), .A2(G146), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n205), .A3(G128), .A4(new_n210), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n208), .A2(new_n211), .B1(new_n194), .B2(new_n193), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT11), .B1(new_n188), .B2(new_n189), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n191), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n188), .B2(new_n189), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(KEYINPUT11), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n213), .B1(new_n218), .B2(new_n187), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G134), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n189), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT11), .B1(new_n223), .B2(new_n215), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n222), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n224), .A2(new_n213), .A3(new_n187), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n195), .B(new_n212), .C1(new_n219), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n215), .B1(new_n226), .B2(G137), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n187), .B(new_n227), .C1(new_n236), .C2(new_n225), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT66), .ZN(new_n238));
  INV_X1    g052(.A(new_n218), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n238), .A2(new_n228), .B1(new_n239), .B2(G131), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n209), .A2(G128), .A3(new_n210), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT0), .ZN(new_n242));
  INV_X1    g056(.A(new_n204), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G128), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n230), .B(new_n235), .C1(new_n240), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G237), .ZN(new_n247));
  INV_X1    g061(.A(G953), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G210), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n249), .B(G101), .Z(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n251));
  XOR2_X1   g065(.A(new_n250), .B(new_n251), .Z(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n238), .A2(new_n228), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n256), .A2(new_n195), .A3(new_n212), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n239), .A2(G131), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n245), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n235), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n230), .B(KEYINPUT30), .C1(new_n240), .C2(new_n245), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n246), .A2(new_n264), .A3(new_n252), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n254), .A2(new_n263), .A3(new_n269), .A4(new_n265), .ZN(new_n270));
  INV_X1    g084(.A(new_n252), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n261), .B1(new_n257), .B2(new_n259), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n246), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n246), .A2(new_n272), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n266), .A2(new_n278), .A3(KEYINPUT31), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n268), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n268), .A2(new_n277), .A3(KEYINPUT71), .A4(new_n279), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n282), .A2(new_n287), .A3(new_n283), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n274), .A2(new_n275), .A3(new_n271), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n295), .B2(KEYINPUT29), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n296), .A2(KEYINPUT75), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n263), .A2(new_n246), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT74), .B1(new_n301), .B2(new_n271), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n299), .B(new_n300), .C1(new_n295), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(KEYINPUT75), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G472), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT76), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .A4(new_n284), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n309), .A3(G472), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n292), .A2(new_n294), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n292), .A2(new_n315), .A3(new_n294), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n319), .A2(KEYINPUT79), .A3(KEYINPUT16), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT79), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n320), .B(new_n321), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(new_n199), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n207), .A2(G119), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(KEYINPUT78), .B2(KEYINPUT23), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n207), .A2(G119), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n329), .A2(new_n332), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n326), .A2(new_n199), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n341));
  INV_X1    g155(.A(new_n203), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n325), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT22), .B(G137), .ZN(new_n345));
  INV_X1    g159(.A(G221), .ZN(new_n346));
  INV_X1    g160(.A(G234), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n346), .A2(new_n347), .A3(G953), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n345), .B(new_n348), .Z(new_n349));
  XNOR2_X1  g163(.A(new_n344), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(KEYINPUT25), .Z(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(G217), .C1(new_n347), .C2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT80), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n347), .B2(G217), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  XNOR2_X1  g176(.A(G110), .B(G122), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT85), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(KEYINPUT82), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(G107), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n368), .B(new_n369), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n371), .A2(G101), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(G101), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n261), .ZN(new_n376));
  INV_X1    g190(.A(new_n369), .ZN(new_n377));
  OAI21_X1  g191(.A(G101), .B1(new_n377), .B2(new_n366), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n378), .A2(KEYINPUT83), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n231), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(new_n233), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G113), .ZN(new_n387));
  INV_X1    g201(.A(G116), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G119), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n376), .B1(KEYINPUT84), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n392), .A2(KEYINPUT84), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n364), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(new_n364), .C1(new_n393), .C2(new_n394), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n393), .A2(new_n394), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n363), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n397), .B(new_n399), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n245), .A2(G125), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n208), .A2(new_n323), .A3(new_n211), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n248), .A2(G224), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n406), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n407), .A2(KEYINPUT7), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n405), .A2(KEYINPUT89), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n413), .B(new_n415), .C1(new_n412), .C2(KEYINPUT89), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n386), .A2(KEYINPUT87), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n390), .B1(new_n386), .B2(KEYINPUT87), .ZN(new_n418));
  OAI221_X1 g232(.A(new_n381), .B1(new_n382), .B2(new_n233), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  OR3_X1    g233(.A1(new_n381), .A2(KEYINPUT88), .A3(new_n391), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT88), .B1(new_n381), .B2(new_n391), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n363), .B(KEYINPUT8), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n414), .B(new_n416), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n424), .B2(new_n401), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n410), .A2(new_n411), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n411), .B1(new_n410), .B2(new_n425), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT90), .B(new_n362), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n425), .ZN(new_n431));
  INV_X1    g245(.A(new_n411), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n426), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT90), .B1(new_n434), .B2(new_n362), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G952), .ZN(new_n437));
  AOI211_X1 g251(.A(G953), .B(new_n437), .C1(G234), .C2(G237), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n351), .B(new_n248), .C1(G234), .C2(G237), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(KEYINPUT95), .B2(KEYINPUT20), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n247), .A2(new_n248), .A3(G214), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n196), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n325), .B(KEYINPUT91), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(G146), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n342), .A2(new_n325), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n326), .A2(new_n199), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n448), .B(G131), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n455), .B(new_n340), .C1(new_n456), .C2(KEYINPUT17), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(KEYINPUT17), .A3(G131), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT93), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n454), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n365), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n451), .A2(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT19), .B2(new_n325), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n467), .A2(new_n468), .A3(new_n342), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n467), .B2(new_n342), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n340), .A3(new_n456), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n462), .B1(new_n471), .B2(new_n454), .ZN(new_n472));
  OAI221_X1 g286(.A(new_n446), .B1(KEYINPUT95), .B2(new_n445), .C1(new_n465), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n445), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n465), .A2(new_n472), .A3(KEYINPUT94), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT94), .B1(new_n465), .B2(new_n472), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G475), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n460), .B(new_n463), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n351), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n479), .A2(KEYINPUT96), .A3(new_n483), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n388), .A2(G122), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT98), .Z(new_n492));
  NOR2_X1   g306(.A1(new_n388), .A2(G122), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n489), .B2(new_n490), .ZN(new_n495));
  OAI21_X1  g309(.A(G107), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G128), .B(G143), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n188), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n226), .A2(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n489), .A2(new_n493), .ZN(new_n502));
  INV_X1    g316(.A(G107), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n502), .B(new_n503), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT97), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT13), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n196), .A3(G128), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n498), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n500), .B1(new_n510), .B2(new_n191), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n505), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT9), .B(G234), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(G217), .A3(new_n248), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n512), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n351), .ZN(new_n516));
  INV_X1    g330(.A(G478), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n516), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n488), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n245), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n375), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n208), .A2(new_n211), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n240), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n209), .A2(new_n210), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n207), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n211), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT10), .B1(new_n381), .B2(new_n529), .ZN(new_n530));
  OR3_X1    g344(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G140), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n248), .A2(G227), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n381), .A2(new_n529), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n523), .B2(new_n381), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n526), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT12), .Z(new_n539));
  AND2_X1   g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n526), .B1(new_n525), .B2(new_n530), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n351), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n351), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n541), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n539), .A2(new_n531), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n546), .B(new_n548), .C1(new_n545), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n346), .B1(new_n513), .B2(new_n351), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n444), .A2(new_n520), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n317), .A2(new_n361), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G101), .ZN(G3));
  NAND3_X1  g372(.A1(new_n282), .A2(new_n351), .A3(new_n284), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G472), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n289), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n360), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n434), .A2(new_n362), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n443), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n515), .A2(new_n517), .A3(new_n351), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n517), .A2(new_n351), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n514), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n515), .B(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n566), .B(new_n568), .C1(new_n572), .C2(new_n517), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n486), .B2(new_n487), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n562), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT34), .B(G104), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  NOR2_X1   g393(.A1(new_n477), .A2(new_n478), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n477), .A2(new_n478), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n482), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n519), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n565), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n562), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G107), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G9));
  INV_X1    g403(.A(new_n349), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n344), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n356), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n355), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n556), .A2(new_n289), .A3(new_n560), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G110), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n595), .B(new_n597), .ZN(G12));
  INV_X1    g412(.A(new_n555), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n564), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT101), .B(G900), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n438), .B1(new_n440), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n585), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n317), .A2(new_n594), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G128), .ZN(G30));
  XOR2_X1   g420(.A(new_n603), .B(KEYINPUT39), .Z(new_n607));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT40), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n293), .B1(new_n289), .B2(new_n290), .ZN(new_n610));
  AOI211_X1 g424(.A(KEYINPUT73), .B(KEYINPUT32), .C1(new_n286), .C2(new_n288), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n266), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n273), .A2(new_n246), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n271), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n616), .B2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(new_n308), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n434), .B(KEYINPUT38), .Z(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n594), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n488), .A2(new_n519), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n362), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n619), .A2(new_n620), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n609), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n196), .ZN(G45));
  INV_X1    g445(.A(new_n603), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n574), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT104), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n317), .A2(new_n594), .A3(new_n601), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G146), .ZN(G48));
  AOI21_X1  g450(.A(new_n360), .B1(new_n314), .B2(new_n316), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n545), .A2(KEYINPUT105), .ZN(new_n638));
  OR3_X1    g452(.A1(new_n543), .A2(G902), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(new_n543), .B2(G902), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n639), .A2(new_n554), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n576), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT41), .B(G113), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G15));
  NAND3_X1  g458(.A1(new_n637), .A2(new_n586), .A3(new_n641), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT106), .B(G116), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G18));
  INV_X1    g461(.A(new_n594), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n314), .B2(new_n316), .ZN(new_n649));
  INV_X1    g463(.A(new_n520), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT107), .B1(new_n641), .B2(new_n564), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n639), .A2(new_n554), .A3(new_n640), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n563), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n649), .A2(new_n443), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  NAND2_X1  g471(.A1(new_n277), .A2(new_n267), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n283), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT108), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(G472), .B2(new_n559), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n358), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n565), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n623), .A4(new_n641), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G122), .ZN(G24));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n594), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT109), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n634), .A3(new_n655), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G125), .ZN(G27));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n555), .B(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n434), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n362), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n634), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n637), .A2(new_n672), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n285), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n312), .B1(new_n679), .B2(KEYINPUT32), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n358), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n672), .A2(new_n681), .A3(new_n634), .A4(new_n675), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n670), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n637), .A2(new_n672), .A3(new_n675), .ZN(new_n686));
  INV_X1    g500(.A(new_n677), .ZN(new_n687));
  OAI211_X1 g501(.A(KEYINPUT111), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G131), .ZN(G33));
  NAND4_X1  g504(.A1(new_n637), .A2(new_n604), .A3(new_n672), .A4(new_n675), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G134), .ZN(G36));
  INV_X1    g506(.A(new_n573), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n488), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n561), .A3(new_n594), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n675), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n551), .B(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G469), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT46), .A3(new_n548), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n546), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT46), .B1(new_n701), .B2(new_n548), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n554), .B(new_n607), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n189), .ZN(G39));
  OAI21_X1  g521(.A(new_n554), .B1(new_n703), .B2(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT47), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n314), .A2(new_n316), .A3(new_n634), .A4(new_n675), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n361), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n318), .ZN(G42));
  INV_X1    g526(.A(new_n694), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n358), .A3(new_n362), .A4(new_n554), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n619), .A2(new_n620), .B1(KEYINPUT112), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n639), .A2(new_n640), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT49), .Z(new_n717));
  OR2_X1    g531(.A1(new_n714), .A2(KEYINPUT112), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n621), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n619), .A2(new_n620), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n674), .A2(new_n652), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n361), .A3(new_n438), .A4(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT116), .Z(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n488), .A3(new_n573), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n696), .A2(new_n438), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n662), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n652), .A2(new_n362), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT115), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n726), .A2(new_n621), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n729), .A2(KEYINPUT50), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(KEYINPUT50), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n725), .A2(new_n721), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n730), .A2(new_n731), .B1(new_n667), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n709), .B1(new_n554), .B2(new_n716), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT117), .Z(new_n735));
  AND2_X1   g549(.A1(new_n726), .A2(new_n675), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n437), .B(G953), .C1(new_n723), .C2(new_n574), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n668), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n648), .B(new_n600), .C1(new_n314), .C2(new_n316), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n634), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n624), .A2(new_n673), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n594), .A2(new_n603), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n618), .A2(new_n744), .A3(new_n599), .A4(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(KEYINPUT52), .A3(new_n605), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n605), .A2(new_n635), .A3(new_n668), .A4(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n656), .A2(new_n642), .A3(new_n645), .A4(new_n664), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT90), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n563), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n574), .A3(new_n443), .A4(new_n429), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n436), .A2(KEYINPUT113), .A3(new_n443), .A4(new_n574), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n488), .A2(new_n584), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n758), .B(new_n759), .C1(new_n444), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n562), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n691), .A2(new_n557), .A3(new_n595), .A4(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n583), .A2(new_n519), .A3(new_n632), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n649), .A2(new_n599), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n672), .A2(new_n667), .A3(new_n634), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n674), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n751), .A2(new_n689), .A3(new_n753), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT54), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n726), .A2(new_n655), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n770), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n315), .B1(new_n612), .B2(new_n312), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT77), .A4(new_n311), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n594), .B(new_n764), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n766), .B1(new_n778), .B2(new_n555), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n675), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n557), .A2(new_n762), .A3(new_n595), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n691), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n750), .B2(new_n747), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n678), .A2(new_n683), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n784), .A4(new_n753), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n775), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n740), .A2(new_n773), .A3(new_n774), .A4(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n724), .A2(new_n733), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n736), .A2(new_n734), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n732), .A2(new_n681), .ZN(new_n793));
  XNOR2_X1  g607(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n789), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(G952), .A2(G953), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n719), .B1(new_n796), .B2(new_n797), .ZN(G75));
  NAND2_X1  g612(.A1(new_n437), .A2(G953), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT120), .Z(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n403), .B(new_n409), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT55), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n351), .B1(new_n775), .B2(new_n785), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(G210), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n805), .B2(KEYINPUT119), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n805), .B(new_n807), .C1(KEYINPUT119), .C2(new_n803), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n801), .B1(new_n809), .B2(new_n810), .ZN(G51));
  AOI211_X1 g625(.A(new_n351), .B(new_n701), .C1(new_n775), .C2(new_n785), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n547), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n775), .A2(new_n785), .A3(new_n787), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n787), .B1(new_n775), .B2(new_n785), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n812), .B1(new_n817), .B2(new_n544), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT122), .B1(new_n818), .B2(new_n801), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n751), .A2(KEYINPUT53), .A3(new_n784), .A4(new_n768), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n752), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n786), .B1(new_n771), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n788), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n543), .B1(new_n824), .B2(new_n814), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n820), .B(new_n800), .C1(new_n825), .C2(new_n812), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n826), .ZN(G54));
  NAND2_X1  g641(.A1(new_n775), .A2(new_n785), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n475), .A2(new_n476), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n804), .A2(KEYINPUT58), .A3(G475), .A4(new_n830), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n800), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(G60));
  XNOR2_X1  g650(.A(new_n567), .B(KEYINPUT59), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n824), .A2(new_n572), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n773), .B2(new_n788), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n839), .B(new_n800), .C1(new_n572), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(G63));
  NAND2_X1  g656(.A1(G217), .A2(G902), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT60), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n775), .B2(new_n785), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n801), .B1(new_n845), .B2(new_n592), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n350), .B2(new_n845), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(G66));
  NAND2_X1  g663(.A1(new_n442), .A2(G224), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(G953), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n753), .A2(new_n781), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(G953), .ZN(new_n853));
  INV_X1    g667(.A(new_n403), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(G898), .B2(new_n248), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n853), .B(new_n855), .ZN(G69));
  NAND2_X1  g670(.A1(new_n260), .A2(new_n262), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(new_n467), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n605), .A2(new_n635), .A3(new_n668), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n861), .C1(new_n630), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n609), .ZN(new_n865));
  INV_X1    g679(.A(new_n629), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n626), .A2(new_n627), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  NAND2_X1  g683(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n862), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n711), .ZN(new_n873));
  INV_X1    g687(.A(new_n608), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n637), .A2(new_n675), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n575), .B2(new_n760), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n706), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(KEYINPUT125), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n711), .B1(new_n864), .B2(new_n871), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n877), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n248), .B(new_n859), .C1(new_n879), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n681), .A2(new_n744), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n705), .B1(new_n699), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n873), .A2(new_n862), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n689), .A2(new_n691), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT126), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n689), .A4(new_n691), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n248), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n858), .C1(G900), .C2(new_n248), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n883), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n248), .B1(G227), .B2(G900), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n883), .A2(new_n895), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(G72));
  NAND3_X1  g715(.A1(new_n889), .A2(new_n852), .A3(new_n892), .ZN(new_n902));
  NAND2_X1  g716(.A1(G472), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT63), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n301), .B(KEYINPUT127), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n271), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n301), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n266), .B1(new_n908), .B2(new_n252), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n904), .B(new_n909), .C1(new_n771), .C2(new_n772), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n800), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n882), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n881), .A2(new_n880), .A3(new_n877), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n852), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n914), .B2(new_n904), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n252), .ZN(G57));
endmodule


