//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n438, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G132), .A4(new_n438), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(G2104), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g040(.A(G101), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n470), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n479), .B2(new_n480), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n490), .B2(new_n495), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n463), .A3(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n481), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n501), .A2(new_n463), .A3(G138), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n469), .A2(new_n504), .A3(KEYINPUT69), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n463), .C1(new_n479), .C2(new_n480), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n505), .B1(KEYINPUT4), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n499), .A2(new_n507), .A3(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n481), .A2(new_n500), .A3(new_n502), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n469), .B2(new_n504), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n488), .B1(new_n467), .B2(new_n468), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n463), .A2(G114), .ZN(new_n515));
  OAI21_X1  g090(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT68), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n509), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n508), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(G164));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT71), .B1(new_n524), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(G543), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G50), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n531), .A2(new_n535), .ZN(new_n538));
  INV_X1    g113(.A(G88), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n534), .A2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND3_X1  g117(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n536), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g121(.A(G89), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n543), .B(new_n544), .C1(new_n548), .C2(KEYINPUT72), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(KEYINPUT72), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(G168));
  AOI22_X1  g126(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n536), .A2(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n538), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n553), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  AOI22_X1  g133(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n533), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n536), .A2(G43), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n538), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  XNOR2_X1  g144(.A(KEYINPUT73), .B(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n531), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(G651), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n536), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OR3_X1    g154(.A1(new_n578), .A2(KEYINPUT9), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  INV_X1    g156(.A(new_n538), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n580), .A2(new_n581), .B1(G91), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n582), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n536), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n536), .A2(G48), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n529), .A2(G86), .A3(new_n530), .A4(new_n535), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n529), .A2(G61), .A3(new_n530), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT75), .Z(new_n595));
  AOI21_X1  g170(.A(new_n533), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n533), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n536), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n538), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n582), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n538), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n536), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT76), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n531), .B2(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n612), .B1(new_n615), .B2(new_n533), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n606), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n606), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(G868), .B2(new_n625), .ZN(G280));
  XOR2_X1   g201(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n564), .B2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n621), .A2(new_n628), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  MUX2_X1   g207(.A(KEYINPUT79), .B(new_n630), .S(new_n632), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g209(.A1(new_n464), .A2(new_n465), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n469), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n477), .A2(G135), .B1(new_n482), .B2(G123), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n645), .A2(new_n463), .A3(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n463), .B2(G111), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT84), .B(G2096), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n642), .A2(new_n643), .A3(new_n651), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2084), .B(G2090), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G2072), .A2(G2078), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n444), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2096), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT20), .Z(new_n691));
  OR2_X1    g266(.A1(new_n684), .A2(new_n686), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(new_n689), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n691), .B1(new_n692), .B2(new_n689), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n697), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n701), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n702), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n702), .B2(new_n706), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(G23), .ZN(new_n718));
  INV_X1    g293(.A(G288), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n714), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT33), .B(G1976), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G6), .A2(G16), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n597), .B2(G16), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n717), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n714), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n604), .B2(new_n714), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(new_n708), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G119), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n738));
  INV_X1    g313(.A(G131), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n738), .C1(new_n739), .C2(new_n470), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n735), .B1(new_n745), .B2(new_n734), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n729), .A2(new_n730), .A3(new_n733), .A4(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT36), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n714), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n714), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n734), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n734), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  OAI21_X1  g333(.A(G29), .B1(new_n472), .B2(new_n475), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n734), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT97), .B(G28), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(KEYINPUT30), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n765), .B2(KEYINPUT30), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n649), .C2(new_n734), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n757), .A2(new_n764), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n734), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT28), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n482), .A2(G128), .ZN(new_n775));
  INV_X1    g350(.A(G140), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n463), .A2(G116), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n775), .B1(new_n776), .B2(new_n470), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT94), .B(G2067), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n759), .A2(new_n763), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2084), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT26), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G129), .B2(new_n482), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n477), .A2(G141), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n635), .A2(G105), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n734), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n734), .B2(G32), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n793), .A2(new_n794), .B1(new_n780), .B2(new_n781), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n753), .A2(new_n772), .A3(new_n784), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G19), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n797), .A2(KEYINPUT93), .A3(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT93), .B1(new_n797), .B2(G16), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(new_n564), .C2(new_n714), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  NOR2_X1   g376(.A1(G27), .A2(G29), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G164), .B2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G2078), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n793), .A2(new_n794), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n734), .A2(G33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n469), .A2(G127), .ZN(new_n808));
  NAND2_X1  g383(.A1(G115), .A2(G2104), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n463), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT25), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n477), .A2(G139), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(KEYINPUT95), .B2(new_n810), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n807), .B1(new_n816), .B2(new_n734), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G2072), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n796), .A2(new_n801), .A3(new_n804), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n714), .A2(G4), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n621), .B2(new_n714), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n714), .A2(G20), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT23), .Z(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G299), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1956), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n714), .A2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G168), .B2(new_n714), .ZN(new_n830));
  INV_X1    g405(.A(G1966), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n824), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n750), .A2(new_n820), .A3(new_n833), .ZN(G311));
  INV_X1    g409(.A(G311), .ZN(G150));
  NOR2_X1   g410(.A1(new_n620), .A2(new_n628), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n560), .A2(new_n563), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n533), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n536), .A2(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n538), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n840), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(G860), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n846), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n851), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(G145));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n779), .B(new_n790), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n514), .A2(new_n517), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n513), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n816), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n816), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n744), .B(new_n638), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n477), .A2(G142), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n463), .A2(KEYINPUT102), .A3(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT102), .B1(new_n463), .B2(G118), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n868), .A2(G2104), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n482), .A2(G130), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n866), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n865), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n486), .B(G160), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n649), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n864), .B2(new_n874), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n857), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n878), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n864), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n865), .A3(new_n878), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g467(.A(new_n631), .B(new_n847), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n621), .A2(G299), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n620), .A2(new_n625), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n894), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n904), .B2(new_n893), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n719), .B(G303), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n604), .B(G305), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n897), .B(new_n909), .C1(new_n904), .C2(new_n893), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G868), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(G868), .B2(new_n853), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  XNOR2_X1  g491(.A(G331), .B(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n847), .A2(G171), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n846), .B(new_n564), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G301), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n920), .A3(G168), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G286), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n902), .A2(new_n903), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n908), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  AOI21_X1  g501(.A(G168), .B1(new_n918), .B2(new_n920), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n894), .B(new_n895), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n857), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n925), .B1(new_n924), .B2(new_n928), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT43), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n935), .A2(new_n894), .A3(new_n895), .ZN(new_n936));
  INV_X1    g511(.A(new_n900), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n925), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n857), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n939), .A2(new_n932), .A3(KEYINPUT43), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n930), .B2(new_n932), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n945), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g521(.A(G1384), .B1(new_n513), .B2(new_n859), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT45), .ZN(new_n948));
  INV_X1    g523(.A(G40), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n472), .A2(new_n475), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n779), .B(G2067), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT107), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n790), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n744), .B(new_n747), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n604), .A2(new_n708), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n951), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT48), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n951), .B1(new_n953), .B2(new_n791), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT124), .ZN(new_n965));
  INV_X1    g540(.A(new_n951), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n954), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT47), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n747), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n956), .A2(new_n971), .B1(G2067), .B2(new_n779), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n963), .B(new_n970), .C1(new_n966), .C2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n604), .A2(new_n708), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n975), .A2(KEYINPUT106), .A3(new_n960), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n966), .B1(new_n975), .B2(KEYINPUT106), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n959), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n950), .B1(new_n947), .B2(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT70), .B1(new_n499), .B2(new_n507), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n513), .A2(new_n520), .A3(new_n509), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(KEYINPUT45), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n985), .B2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n522), .A2(new_n987), .A3(KEYINPUT45), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n831), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(new_n859), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n983), .B1(new_n507), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n950), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n992), .A2(new_n758), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(G168), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1966), .B1(new_n986), .B2(new_n988), .ZN(new_n1000));
  OAI21_X1  g575(.A(G286), .B1(new_n1000), .B2(new_n997), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(G8), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT51), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1004), .A3(G8), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n719), .A2(G1976), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n947), .A2(new_n950), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(KEYINPUT109), .A3(G8), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT109), .B1(new_n1012), .B2(G8), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1009), .B(new_n1011), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n593), .A2(new_n595), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G651), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(new_n703), .A3(new_n591), .A4(new_n590), .ZN(new_n1019));
  OAI21_X1  g594(.A(G1981), .B1(new_n592), .B2(new_n596), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1014), .A2(new_n1015), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1012), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1013), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1030), .B2(new_n1009), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n992), .A2(new_n996), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2090), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n950), .B1(new_n994), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1040), .B2(new_n991), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT108), .B(G1971), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1037), .B(G8), .C1(new_n1039), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1032), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n982), .A2(new_n1047), .A3(new_n983), .A4(new_n984), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n473), .A2(new_n474), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G2105), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n477), .A2(G137), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(G40), .A4(new_n466), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1042), .A2(new_n1043), .B1(new_n1054), .B2(G2090), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1037), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1008), .B1(new_n1046), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n995), .B1(KEYINPUT50), .B2(new_n991), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G1961), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n991), .A2(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1041), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G2078), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n986), .A2(new_n988), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(G301), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1032), .A2(new_n1058), .A3(KEYINPUT121), .A4(new_n1045), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1060), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1007), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1045), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1032), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n719), .A2(new_n1010), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1030), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1019), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1030), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1083), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1079), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1032), .A2(new_n1045), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT112), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(G8), .C1(new_n1039), .C2(new_n1044), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1057), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G168), .A2(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n990), .B2(new_n998), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(new_n1094), .A3(KEYINPUT63), .A4(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1032), .A2(new_n1096), .A3(new_n1058), .A4(new_n1045), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1088), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1063), .A2(new_n1064), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT115), .B1(new_n1042), .B2(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT113), .B(G1956), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1054), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT114), .B(new_n1108), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1105), .A2(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n577), .A2(new_n583), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n577), .B2(new_n583), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  OAI221_X1 g695(.A(new_n1117), .B1(new_n1110), .B2(new_n1111), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1042), .A2(KEYINPUT115), .A3(new_n1102), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1054), .A2(new_n1109), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1054), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1123), .A2(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT117), .B(G1996), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1042), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1012), .A2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n1131), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1065), .B2(new_n1132), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1131), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1012), .ZN(new_n1143));
  INV_X1    g718(.A(G2067), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT60), .B(new_n1145), .C1(new_n1061), .C2(G1348), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(KEYINPUT119), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(KEYINPUT119), .A3(new_n620), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n620), .B1(new_n1146), .B2(KEYINPUT119), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1145), .B1(new_n1061), .B2(G1348), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1142), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT116), .B1(new_n1128), .B2(new_n1117), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1112), .A2(new_n1118), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1151), .A2(new_n621), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1130), .A2(new_n1154), .B1(new_n1159), .B2(new_n1121), .ZN(new_n1160));
  OAI221_X1 g735(.A(new_n1071), .B1(G1961), .B2(new_n1061), .C1(new_n1066), .C2(KEYINPUT53), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G301), .B(KEYINPUT54), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1070), .B1(new_n994), .B2(new_n1040), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n981), .A2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1165), .A2(new_n1166), .A3(new_n1162), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1161), .A2(new_n1162), .B1(new_n1069), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1006), .A2(new_n1060), .A3(new_n1073), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1101), .B1(new_n1160), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1077), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1101), .B(KEYINPUT122), .C1(new_n1160), .C2(new_n1169), .ZN(new_n1173));
  AOI211_X1 g748(.A(KEYINPUT123), .B(new_n980), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1077), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n1173), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n979), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n973), .B1(new_n1174), .B2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n1182));
  OAI21_X1  g756(.A(G319), .B1(new_n666), .B2(new_n667), .ZN(new_n1183));
  NOR2_X1   g757(.A1(G227), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g758(.A(new_n1184), .B(KEYINPUT125), .Z(new_n1185));
  OAI211_X1 g759(.A(new_n712), .B(new_n1185), .C1(new_n889), .C2(new_n884), .ZN(new_n1186));
  AOI211_X1 g760(.A(new_n1182), .B(new_n1186), .C1(new_n943), .C2(new_n944), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n944), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1186), .ZN(new_n1189));
  AOI21_X1  g763(.A(KEYINPUT126), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1187), .A2(new_n1190), .ZN(G308));
  OAI21_X1  g765(.A(new_n1182), .B1(new_n945), .B2(new_n1186), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n1188), .A2(KEYINPUT126), .A3(new_n1189), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1193), .ZN(G225));
endmodule


