//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT77), .A2(G101), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT77), .A2(G101), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n188), .A2(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(new_n192), .A3(new_n198), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(new_n196), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT78), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n191), .A2(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n199), .A2(new_n202), .B1(G101), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(G128), .B1(new_n213), .B2(new_n208), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n212), .A2(G143), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(KEYINPUT66), .C1(G128), .C2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n220), .B(G128), .C1(new_n210), .C2(new_n209), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OR3_X1    g037(.A1(new_n205), .A2(KEYINPUT79), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n222), .B(new_n225), .C1(G128), .C2(new_n220), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n205), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT79), .B1(new_n205), .B2(new_n223), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n200), .A2(G101), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n199), .A2(new_n202), .B1(G101), .B2(new_n200), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n242), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  AND2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  OR3_X1    g062(.A1(new_n220), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n237), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n227), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n205), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n250), .A2(new_n251), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n229), .A2(new_n237), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n240), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n259), .B(new_n261), .Z(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n255), .A2(new_n262), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n237), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G469), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n257), .ZN(new_n272));
  INV_X1    g086(.A(new_n239), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n229), .B2(new_n237), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT82), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n240), .A2(new_n276), .A3(new_n257), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n277), .A3(new_n265), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n255), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n263), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n270), .A3(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n258), .A2(new_n263), .B1(new_n267), .B2(new_n265), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT81), .B(G469), .C1(new_n284), .C2(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n271), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT9), .B(G234), .Z(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G221), .B1(new_n288), .B2(G902), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G475), .ZN(new_n291));
  XNOR2_X1  g105(.A(G125), .B(G140), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT16), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  OR3_X1    g108(.A1(new_n294), .A2(KEYINPUT16), .A3(G140), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(G146), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G146), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G237), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n260), .A3(G214), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(G143), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT17), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n302), .B(new_n303), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n299), .B(new_n305), .C1(new_n306), .C2(KEYINPUT17), .ZN(new_n307));
  XNOR2_X1  g121(.A(G113), .B(G122), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(new_n188), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(KEYINPUT18), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT18), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n302), .B1(new_n311), .B2(new_n303), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n292), .B(new_n212), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n307), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n292), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT19), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n292), .A2(new_n317), .A3(KEYINPUT19), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n316), .B(new_n296), .C1(new_n322), .C2(G146), .ZN(new_n323));
  AOI21_X1  g137(.A(G146), .B1(new_n320), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT89), .B1(new_n324), .B2(new_n297), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(new_n306), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n309), .B1(new_n326), .B2(new_n314), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n291), .B(new_n282), .C1(new_n315), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT20), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT90), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT20), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n328), .A2(KEYINPUT20), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n309), .B1(new_n307), .B2(new_n314), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n282), .B1(new_n315), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G475), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G128), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G143), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n207), .A2(G128), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n231), .ZN(new_n343));
  XNOR2_X1  g157(.A(G116), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n191), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT13), .B1(new_n207), .B2(G128), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n341), .B(new_n348), .C1(KEYINPUT13), .C2(new_n340), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n343), .B(new_n345), .C1(new_n349), .C2(new_n231), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n342), .B(new_n231), .ZN(new_n351));
  INV_X1    g165(.A(G116), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT14), .A3(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n344), .ZN(new_n354));
  OAI211_X1 g168(.A(G107), .B(new_n353), .C1(new_n354), .C2(KEYINPUT14), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n351), .B(new_n355), .C1(G107), .C2(new_n354), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n288), .A2(new_n358), .A3(G953), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n350), .A2(new_n356), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n282), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT93), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n364), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(KEYINPUT93), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n364), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n260), .A2(G952), .ZN(new_n374));
  NAND2_X1  g188(.A1(G234), .A2(G237), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT21), .B(G898), .Z(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(G902), .A3(G953), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n338), .A2(new_n373), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(G110), .B(G122), .Z(new_n384));
  INV_X1    g198(.A(G119), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G116), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n352), .A2(G119), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n389));
  XNOR2_X1  g203(.A(G116), .B(G119), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT69), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT5), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n394));
  INV_X1    g208(.A(G113), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT68), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT2), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n399), .A2(new_n400), .B1(KEYINPUT2), .B2(G113), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n393), .A2(new_n396), .B1(new_n401), .B2(new_n390), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n390), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n389), .A2(new_n392), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n401), .ZN(new_n405));
  AOI221_X4 g219(.A(KEYINPUT83), .B1(new_n205), .B2(new_n402), .C1(new_n245), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n199), .A2(new_n202), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n242), .B1(new_n408), .B2(new_n241), .ZN(new_n409));
  INV_X1    g223(.A(new_n243), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n205), .A2(new_n402), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT6), .B(new_n384), .C1(new_n406), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n384), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n189), .A2(new_n192), .A3(new_n198), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n194), .B1(new_n416), .B2(new_n197), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n200), .A2(KEYINPUT78), .A3(new_n201), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n241), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n410), .B1(new_n419), .B2(KEYINPUT4), .ZN(new_n420));
  INV_X1    g234(.A(new_n405), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n412), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n411), .A2(new_n407), .A3(new_n412), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n245), .A2(new_n405), .B1(new_n205), .B2(new_n402), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n415), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n414), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n260), .A2(G224), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT85), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n223), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n249), .A2(new_n246), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G125), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(G125), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n433), .A2(new_n439), .A3(new_n431), .A4(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n429), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n431), .A2(KEYINPUT7), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n433), .B2(new_n438), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n437), .A2(new_n440), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n427), .A2(new_n415), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n205), .A2(new_n402), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n454));
  INV_X1    g268(.A(new_n396), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n205), .B(new_n403), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n384), .B(KEYINPUT8), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n450), .B(new_n451), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n282), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n429), .A2(new_n443), .A3(KEYINPUT86), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n446), .A2(new_n465), .A3(new_n462), .A4(new_n463), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n383), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n290), .A2(new_n381), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n236), .A2(G131), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n234), .A2(G134), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n303), .B1(new_n233), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT64), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n223), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n237), .A2(new_n246), .A3(new_n249), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n471), .A4(new_n474), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n475), .A2(KEYINPUT70), .A3(new_n478), .A4(KEYINPUT30), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n487), .A3(new_n405), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n482), .A2(new_n487), .A3(new_n490), .A4(new_n405), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n421), .A2(new_n475), .A3(new_n478), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(G101), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n300), .A2(new_n260), .A3(G210), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n492), .A2(KEYINPUT28), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(KEYINPUT28), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n480), .A2(new_n405), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n496), .A2(KEYINPUT29), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n421), .B1(new_n478), .B2(new_n475), .ZN(new_n510));
  AOI211_X1 g324(.A(new_n509), .B(new_n510), .C1(new_n501), .C2(new_n502), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n508), .B1(new_n511), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(KEYINPUT72), .B(new_n282), .C1(new_n514), .C2(new_n509), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G472), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(G472), .C1(new_n507), .C2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n481), .A2(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n490), .B1(new_n522), .B2(new_n405), .ZN(new_n523));
  AND4_X1   g337(.A1(new_n490), .A2(new_n482), .A3(new_n487), .A4(new_n405), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n492), .A4(new_n496), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n505), .A2(new_n497), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n489), .A2(new_n492), .A3(new_n496), .A4(new_n491), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT31), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n521), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n358), .B1(G234), .B2(new_n282), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n385), .B2(G128), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n339), .A2(KEYINPUT23), .A3(G119), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n539), .B(new_n540), .C1(G119), .C2(new_n339), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G110), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT75), .Z(new_n543));
  XNOR2_X1  g357(.A(G119), .B(G128), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n292), .A2(new_n212), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n296), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n299), .B1(new_n544), .B2(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(G110), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT22), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(G137), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n548), .A2(new_n552), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT25), .B1(new_n561), .B2(new_n282), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n560), .A2(new_n563), .A3(G902), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n537), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n282), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n566), .A2(new_n537), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n536), .A2(KEYINPUT76), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT76), .B1(new_n536), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n470), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n201), .ZN(G3));
  NAND2_X1  g386(.A1(new_n531), .A2(new_n533), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n565), .B1(new_n537), .B2(new_n566), .ZN(new_n575));
  INV_X1    g389(.A(G472), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n531), .B2(new_n282), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n290), .ZN(new_n579));
  INV_X1    g393(.A(new_n338), .ZN(new_n580));
  INV_X1    g394(.A(new_n362), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n359), .B1(new_n350), .B2(new_n356), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT33), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n361), .A2(new_n584), .A3(new_n362), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n585), .A3(G478), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n363), .A2(new_n366), .A3(new_n282), .ZN(new_n587));
  NAND2_X1  g401(.A1(G478), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n469), .A2(new_n379), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n469), .A2(KEYINPUT94), .A3(new_n379), .A4(new_n590), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n579), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT34), .B(G104), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  XOR2_X1   g411(.A(new_n379), .B(KEYINPUT96), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n383), .B(new_n599), .C1(new_n467), .C2(new_n468), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n373), .A2(new_n337), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n333), .B(KEYINPUT95), .Z(new_n602));
  AND2_X1   g416(.A1(new_n330), .A2(new_n332), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n579), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT97), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n606), .B(new_n608), .ZN(G9));
  NAND2_X1  g423(.A1(new_n531), .A2(new_n282), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n553), .B(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n282), .C1(new_n358), .C2(G234), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n565), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n611), .A2(new_n573), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(new_n381), .A3(new_n469), .A4(new_n290), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT98), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT37), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  NAND2_X1  g434(.A1(new_n467), .A2(new_n468), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n382), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n625), .B2(new_n521), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n376), .B1(G900), .B2(new_n378), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n604), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n286), .A2(new_n289), .A3(new_n615), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  INV_X1    g446(.A(new_n443), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n384), .B1(new_n406), .B2(new_n413), .ZN(new_n634));
  INV_X1    g448(.A(new_n428), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n445), .B(new_n633), .C1(new_n636), .C2(new_n414), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT86), .B1(new_n429), .B2(new_n443), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n465), .B1(new_n639), .B2(new_n462), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n637), .A2(new_n638), .A3(new_n466), .A4(new_n461), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n525), .A2(new_n492), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n496), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n282), .B1(new_n498), .B2(new_n510), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n615), .B1(new_n625), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n338), .A2(new_n373), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n627), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n290), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  AND4_X1   g470(.A1(new_n382), .A2(new_n644), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n207), .ZN(G45));
  INV_X1    g472(.A(new_n627), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n659), .B(new_n589), .C1(new_n334), .C2(new_n337), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n382), .B(new_n660), .C1(new_n640), .C2(new_n641), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n469), .A2(KEYINPUT100), .A3(new_n660), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n629), .B1(new_n625), .B2(new_n521), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n212), .ZN(G48));
  NAND2_X1  g485(.A1(new_n593), .A2(new_n594), .ZN(new_n672));
  INV_X1    g486(.A(new_n283), .ZN(new_n673));
  INV_X1    g487(.A(new_n289), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n270), .B1(new_n281), .B2(new_n282), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n536), .A2(new_n568), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n677), .B2(new_n605), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n575), .B1(new_n625), .B2(new_n521), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n469), .A2(new_n598), .A3(new_n604), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(KEYINPUT102), .A4(new_n676), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT103), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n352), .ZN(G18));
  NAND4_X1  g503(.A1(new_n626), .A2(new_n381), .A3(new_n615), .A4(new_n676), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND2_X1  g505(.A1(new_n514), .A2(new_n497), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n527), .A2(new_n530), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n533), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT104), .B1(new_n693), .B2(new_n533), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n611), .B(new_n568), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n676), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n651), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n600), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  OAI211_X1 g514(.A(new_n611), .B(new_n615), .C1(new_n694), .C2(new_n695), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n693), .A2(new_n533), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n533), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n611), .A4(new_n615), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n697), .A2(new_n661), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n284), .B2(G902), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n283), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n674), .A2(new_n383), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n642), .A2(new_n714), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n716), .A2(new_n467), .A3(new_n468), .A4(new_n717), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n684), .A3(new_n660), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n590), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n718), .B2(new_n720), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n627), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n303), .ZN(G33));
  AND3_X1   g543(.A1(new_n721), .A2(new_n684), .A3(new_n628), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n231), .ZN(G36));
  OR2_X1    g545(.A1(new_n284), .A2(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n284), .A2(KEYINPUT45), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT107), .Z(new_n735));
  NOR2_X1   g549(.A1(new_n270), .A2(new_n282), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n283), .B1(new_n737), .B2(KEYINPUT46), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n289), .B(new_n654), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n621), .A2(new_n383), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n589), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n580), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT43), .Z(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(new_n615), .C1(new_n574), .C2(new_n577), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n743), .B1(new_n748), .B2(KEYINPUT44), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n741), .B(new_n749), .C1(KEYINPUT44), .C2(new_n748), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  OAI21_X1  g565(.A(new_n289), .B1(new_n738), .B2(new_n739), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT47), .B(new_n289), .C1(new_n738), .C2(new_n739), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n536), .A2(new_n568), .A3(new_n725), .A4(new_n659), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n742), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  INV_X1    g573(.A(new_n376), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n746), .A2(new_n760), .A3(new_n676), .A4(new_n742), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n709), .B2(new_n702), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT113), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n742), .A2(new_n760), .A3(new_n676), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n625), .A2(new_n649), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n764), .A2(new_n765), .A3(new_n575), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n338), .A3(new_n744), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n696), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n746), .A2(new_n769), .A3(new_n760), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n743), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT110), .Z(new_n772));
  NOR2_X1   g586(.A1(new_n673), .A2(new_n675), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n674), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n772), .B1(new_n756), .B2(new_n775), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n644), .A2(new_n382), .A3(new_n697), .A4(new_n770), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT50), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n768), .B(new_n776), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n536), .A2(new_n568), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n761), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT48), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n770), .A2(new_n622), .A3(new_n697), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n374), .C1(new_n725), .C2(new_n766), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT114), .Z(new_n790));
  INV_X1    g604(.A(new_n774), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n772), .B1(new_n756), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n778), .A2(new_n792), .A3(KEYINPUT51), .A4(new_n768), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n783), .A2(new_n796), .A3(new_n790), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n578), .A2(new_n600), .A3(new_n290), .A4(new_n590), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n601), .B1(new_n603), .B2(new_n333), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n578), .A2(new_n600), .A3(new_n290), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n617), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n802), .B1(new_n617), .B2(new_n801), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n571), .B(new_n799), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n672), .A2(new_n678), .B1(new_n698), .B2(new_n600), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n687), .A3(new_n690), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(new_n687), .A3(new_n809), .A4(new_n690), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n631), .B(new_n712), .C1(new_n668), .C2(new_n669), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n650), .A2(new_n289), .A3(new_n627), .ZN(new_n814));
  INV_X1    g628(.A(new_n716), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n469), .A2(new_n652), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n812), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n661), .A2(new_n662), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT100), .B1(new_n469), .B2(new_n660), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n667), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(KEYINPUT52), .A3(new_n712), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n710), .A2(new_n726), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n373), .B1(new_n602), .B2(new_n603), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n337), .A2(new_n667), .A3(new_n742), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n627), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n730), .B1(new_n724), .B2(new_n727), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n811), .A2(new_n828), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n834), .B1(new_n818), .B2(new_n827), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n805), .A2(new_n807), .A3(new_n837), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  OAI22_X1  g660(.A1(new_n798), .A2(new_n846), .B1(G952), .B2(G953), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n644), .A2(new_n383), .A3(new_n674), .A4(new_n745), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n773), .B(KEYINPUT49), .Z(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n575), .A3(new_n765), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n847), .A2(new_n851), .ZN(G75));
  NOR2_X1   g666(.A1(new_n260), .A2(G952), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n840), .A2(new_n844), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(G210), .A3(G902), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n429), .B(new_n443), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT55), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n856), .A2(KEYINPUT56), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n861), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n858), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(KEYINPUT117), .B(new_n858), .C1(new_n860), .C2(new_n863), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n853), .B(new_n859), .C1(new_n866), .C2(new_n867), .ZN(G51));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n842), .B2(new_n811), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n828), .A2(new_n835), .A3(new_n843), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n282), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n735), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n845), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n736), .B(KEYINPUT57), .Z(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT118), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n881), .B(new_n878), .C1(new_n845), .C2(new_n876), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n875), .B1(new_n883), .B2(new_n281), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n869), .B1(new_n884), .B2(new_n853), .ZN(new_n885));
  INV_X1    g699(.A(new_n853), .ZN(new_n886));
  INV_X1    g700(.A(new_n281), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n880), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT119), .B(new_n886), .C1(new_n888), .C2(new_n875), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(G54));
  NAND3_X1  g704(.A1(new_n873), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n315), .A2(new_n327), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n853), .ZN(G60));
  NAND2_X1  g708(.A1(new_n583), .A2(new_n585), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n588), .B(KEYINPUT59), .Z(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n877), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n839), .B2(new_n845), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n886), .B(new_n898), .C1(new_n899), .C2(new_n895), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT120), .Z(G63));
  XNOR2_X1  g715(.A(new_n613), .B(KEYINPUT123), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n358), .A2(new_n282), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT122), .B1(new_n872), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n854), .A2(new_n909), .A3(new_n905), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n902), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n910), .A3(new_n560), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n886), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT124), .B(new_n902), .C1(new_n908), .C2(new_n911), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT61), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(G66));
  AOI21_X1  g736(.A(new_n260), .B1(new_n377), .B2(G224), .ZN(new_n923));
  INV_X1    g737(.A(new_n811), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n260), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n636), .B(new_n414), .C1(G898), .C2(new_n260), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(G69));
  AOI21_X1  g741(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n758), .A2(new_n750), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n657), .A2(KEYINPUT62), .A3(new_n813), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n657), .B2(new_n813), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n569), .A2(new_n570), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n742), .B1(new_n590), .B2(new_n800), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n933), .A2(new_n655), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT125), .B1(new_n936), .B2(new_n260), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n758), .A2(new_n712), .A3(new_n750), .A4(new_n825), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n741), .A2(new_n684), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n833), .B1(new_n939), .B2(new_n816), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n260), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n522), .B(new_n322), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n260), .A2(G900), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n937), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n936), .A2(new_n260), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n947), .B2(KEYINPUT125), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n929), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n946), .A2(new_n948), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n928), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n953), .B(new_n929), .C1(new_n946), .C2(new_n948), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n950), .A2(new_n952), .A3(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n936), .B2(new_n924), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n853), .B1(new_n958), .B2(new_n647), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n938), .A2(new_n940), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n960), .B2(new_n924), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n525), .A3(new_n499), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n838), .A2(new_n500), .A3(new_n646), .A4(new_n957), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(G57));
endmodule


