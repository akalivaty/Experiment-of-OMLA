//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  AOI21_X1  g002(.A(G8gat), .B1(new_n203), .B2(KEYINPUT93), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n205), .A2(new_n206), .A3(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n204), .B(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT91), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n219), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n214), .A3(new_n217), .ZN(new_n226));
  INV_X1    g025(.A(new_n224), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(KEYINPUT91), .C2(new_n218), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT94), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n228), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(KEYINPUT17), .ZN(new_n234));
  AOI211_X1 g033(.A(KEYINPUT94), .B(new_n230), .C1(new_n225), .C2(new_n228), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n211), .B(new_n231), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n211), .A2(new_n233), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n239), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n211), .B(new_n233), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n237), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT11), .B(G169gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n242), .A2(new_n252), .A3(new_n243), .A4(new_n246), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G141gat), .B(G148gat), .Z(new_n258));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT2), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n259), .A2(new_n263), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n259), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(new_n262), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n258), .B(new_n260), .C1(new_n268), .C2(new_n264), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n273), .A2(KEYINPUT68), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(G120gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G113gat), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G120gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT1), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n274), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n273), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT69), .B(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n277), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(KEYINPUT70), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT4), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n266), .A2(new_n269), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT80), .B1(new_n293), .B2(KEYINPUT3), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(KEYINPUT3), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n282), .B(KEYINPUT81), .C1(new_n288), .C2(new_n289), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n290), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n270), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n292), .A2(new_n301), .A3(new_n302), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n298), .A2(new_n299), .ZN(new_n308));
  MUX2_X1   g107(.A(new_n290), .B(new_n308), .S(new_n293), .Z(new_n309));
  OAI211_X1 g108(.A(new_n307), .B(KEYINPUT5), .C1(new_n309), .C2(new_n302), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n270), .B(KEYINPUT82), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT83), .B1(new_n312), .B2(KEYINPUT4), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n314), .A3(new_n305), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(KEYINPUT4), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n302), .A4(new_n301), .ZN(new_n319));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT0), .ZN(new_n321));
  XNOR2_X1  g120(.A(G57gat), .B(G85gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  AND3_X1   g122(.A1(new_n310), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n310), .B2(new_n319), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT6), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT89), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n326), .A2(new_n327), .B1(KEYINPUT6), .B2(new_n325), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n319), .ZN(new_n329));
  INV_X1    g128(.A(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT6), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n319), .A3(new_n323), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT89), .ZN(new_n335));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT74), .B(G218gat), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n347), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT64), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(KEYINPUT24), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G169gat), .ZN(new_n360));
  INV_X1    g159(.A(G176gat), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n360), .A2(new_n361), .B1(KEYINPUT65), .B2(KEYINPUT25), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n358), .A2(KEYINPUT24), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT27), .B(G183gat), .Z(new_n368));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT66), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n368), .A2(G190gat), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT67), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n372), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(KEYINPUT26), .B2(new_n372), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n369), .A2(KEYINPUT66), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n370), .B(new_n375), .C1(new_n368), .C2(G190gat), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(new_n374), .A3(new_n376), .A4(new_n358), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n379));
  AOI21_X1  g178(.A(new_n352), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n351), .B1(new_n367), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n381), .A2(KEYINPUT77), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n350), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n347), .B(new_n348), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n378), .A2(new_n352), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n386), .A2(KEYINPUT78), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n367), .B2(new_n377), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(KEYINPUT78), .C1(new_n352), .C2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n385), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n339), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT37), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n338), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n382), .A2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n385), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n350), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n392), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT38), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(new_n338), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n392), .B1(new_n397), .B2(new_n385), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n350), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT38), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n393), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n328), .A2(new_n335), .A3(new_n400), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G228gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n379), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n385), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n272), .B1(new_n412), .B2(KEYINPUT3), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n379), .B1(new_n293), .B2(KEYINPUT3), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n350), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n410), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n350), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n270), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n385), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n410), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(G22gat), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G78gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n350), .A2(new_n379), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n311), .B1(new_n431), .B2(new_n421), .ZN(new_n432));
  OAI22_X1  g231(.A1(new_n432), .A2(new_n416), .B1(new_n408), .B2(new_n409), .ZN(new_n433));
  INV_X1    g232(.A(G22gat), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT3), .B1(new_n350), .B2(new_n419), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n410), .B(new_n426), .C1(new_n435), .C2(new_n270), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n429), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n429), .B2(new_n437), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT31), .B(G50gat), .ZN(new_n440));
  INV_X1    g239(.A(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n418), .A2(G22gat), .A3(new_n428), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n434), .B1(new_n433), .B2(new_n436), .ZN(new_n446));
  OAI21_X1  g245(.A(G78gat), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n437), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n317), .A2(new_n301), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453));
  INV_X1    g252(.A(new_n302), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n302), .B(new_n304), .C1(new_n308), .C2(new_n270), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT39), .B1(new_n460), .B2(KEYINPUT88), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(KEYINPUT88), .B2(new_n460), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n463), .A3(new_n323), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n458), .A2(new_n463), .A3(KEYINPUT40), .A4(new_n323), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OR4_X1    g267(.A1(KEYINPUT30), .A2(new_n384), .A3(new_n390), .A4(new_n339), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n401), .A2(new_n391), .A3(KEYINPUT30), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n470), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n331), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n407), .B(new_n450), .C1(new_n468), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n325), .A2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n334), .A2(new_n478), .B1(new_n469), .B2(new_n470), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n443), .B1(new_n438), .B2(new_n439), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n447), .A2(new_n448), .A3(new_n442), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n378), .A2(new_n303), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(new_n409), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n367), .A2(new_n290), .A3(new_n377), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  INV_X1    g291(.A(G15gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n487), .B(KEYINPUT32), .C1(new_n489), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n485), .B1(new_n483), .B2(new_n486), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n483), .A2(new_n486), .ZN(new_n506));
  INV_X1    g305(.A(new_n485), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n503), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n505), .A2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n500), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n510), .A2(KEYINPUT36), .A3(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n511), .A2(new_n500), .A3(KEYINPUT73), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n500), .B(new_n509), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n477), .B1(new_n482), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n334), .A2(new_n478), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n471), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n444), .B2(new_n449), .ZN(new_n522));
  INV_X1    g321(.A(new_n513), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(KEYINPUT73), .B2(new_n510), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n525), .B2(KEYINPUT36), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n526), .A3(KEYINPUT85), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n476), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n328), .A2(new_n335), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n473), .A2(new_n474), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n450), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n480), .A2(new_n479), .A3(new_n515), .A4(new_n481), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n257), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(G57gat), .A2(G64gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT9), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  OR3_X1    g340(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545));
  INV_X1    g344(.A(G71gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n430), .A3(KEYINPUT9), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT96), .B1(new_n537), .B2(new_n538), .ZN(new_n548));
  INV_X1    g347(.A(G57gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  NAND2_X1  g351(.A1(G57gat), .A2(G64gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI221_X4 g353(.A(new_n545), .B1(new_n541), .B2(new_n547), .C1(new_n548), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(new_n541), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT97), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n544), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G127gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n211), .B1(new_n560), .B2(new_n559), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n568));
  INV_X1    g367(.A(G155gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n565), .B(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n572), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n233), .A2(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT94), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n233), .A2(new_n232), .A3(KEYINPUT17), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  OAI21_X1  g383(.A(G92gat), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n582), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT8), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(KEYINPUT98), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(KEYINPUT98), .B2(new_n590), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n588), .B2(new_n592), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT99), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n588), .A2(new_n592), .ZN(new_n599));
  INV_X1    g398(.A(new_n593), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n594), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n230), .B2(new_n229), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n229), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n581), .B2(new_n606), .ZN(new_n616));
  INV_X1    g415(.A(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n615), .B2(new_n618), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n599), .A2(new_n626), .A3(new_n593), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n588), .B(new_n592), .C1(KEYINPUT101), .C2(new_n600), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n559), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n542), .A2(new_n541), .A3(new_n543), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(KEYINPUT9), .B2(new_n539), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT96), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n557), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n545), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n556), .A2(KEYINPUT97), .A3(new_n557), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n631), .B1(new_n639), .B2(new_n602), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n559), .A2(new_n597), .A3(KEYINPUT100), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n630), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n639), .A2(KEYINPUT10), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n604), .B2(new_n598), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n647), .B1(new_n651), .B2(new_n645), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n627), .A3(new_n628), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n631), .A3(new_n602), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT100), .B1(new_n559), .B2(new_n597), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n650), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n639), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(KEYINPUT102), .A3(new_n644), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n646), .A2(new_n652), .A3(new_n655), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n655), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n651), .A2(new_n645), .ZN(new_n666));
  INV_X1    g465(.A(new_n646), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n577), .A2(new_n625), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n536), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n520), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  INV_X1    g473(.A(new_n530), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n676), .A2(G8gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT42), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(KEYINPUT42), .B2(new_n679), .ZN(G1325gat));
  INV_X1    g480(.A(new_n671), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n682), .B2(new_n526), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n671), .A2(new_n493), .A3(new_n525), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n480), .A2(new_n481), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n536), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n670), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  INV_X1    g489(.A(new_n577), .ZN(new_n691));
  INV_X1    g490(.A(new_n625), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(new_n692), .A3(new_n669), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n536), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(G29gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n672), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n621), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n613), .A2(new_n614), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n616), .A2(new_n617), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n622), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT106), .B1(new_n703), .B2(new_n622), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n522), .A2(new_n526), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n468), .A2(new_n475), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n326), .A2(new_n327), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n710), .A2(new_n478), .A3(new_n335), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n400), .A2(new_n406), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n686), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n708), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n532), .A2(new_n534), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n707), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n692), .B1(new_n528), .B2(new_n535), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n574), .A2(KEYINPUT105), .A3(new_n576), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n574), .B2(new_n576), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(new_n257), .A3(new_n669), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n520), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(G36gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n694), .A2(new_n728), .A3(new_n675), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT46), .Z(new_n730));
  OAI21_X1  g529(.A(G36gat), .B1(new_n725), .B2(new_n530), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1329gat));
  NOR3_X1   g531(.A1(new_n725), .A2(new_n495), .A3(new_n526), .ZN(new_n733));
  AOI21_X1  g532(.A(G43gat), .B1(new_n694), .B2(new_n525), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g535(.A(G50gat), .B1(new_n725), .B2(new_n450), .ZN(new_n737));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n687), .A2(new_n738), .A3(new_n693), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g540(.A1(new_n476), .A2(new_n522), .A3(new_n526), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n535), .ZN(new_n743));
  INV_X1    g542(.A(new_n669), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n577), .A2(new_n256), .A3(new_n625), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n672), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g547(.A(new_n746), .B(KEYINPUT107), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n530), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  INV_X1    g554(.A(new_n746), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n546), .B1(new_n756), .B2(new_n516), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n518), .A2(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n750), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n749), .A2(new_n686), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g561(.A1(new_n577), .A2(new_n257), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n692), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n743), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n743), .A2(KEYINPUT51), .A3(new_n764), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n744), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n584), .A3(new_n672), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n763), .A2(new_n744), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n719), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n719), .B2(new_n772), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n773), .A2(new_n774), .A3(new_n520), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n775), .B2(new_n584), .ZN(G1336gat));
  NAND2_X1  g575(.A1(new_n719), .A2(new_n772), .ZN(new_n777));
  OAI21_X1  g576(.A(G92gat), .B1(new_n777), .B2(new_n530), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n530), .A2(G92gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n769), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n774), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n719), .A2(new_n771), .A3(new_n772), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n675), .A3(new_n784), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n785), .A2(G92gat), .B1(new_n769), .B2(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n786), .B2(new_n779), .ZN(G1337gat));
  INV_X1    g586(.A(G99gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n788), .A3(new_n525), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n526), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n789), .C1(new_n790), .C2(new_n788), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1338gat));
  OAI21_X1  g594(.A(G106gat), .B1(new_n777), .B2(new_n450), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n450), .A2(G106gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n769), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n686), .A3(new_n784), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(G106gat), .B1(new_n769), .B2(new_n798), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n797), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n623), .B2(new_n624), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n622), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n661), .A2(new_n644), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n665), .B1(new_n808), .B2(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT102), .B1(new_n661), .B2(new_n644), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n647), .B(new_n645), .C1(new_n659), .C2(new_n660), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n651), .B2(new_n645), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n809), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n663), .B1(new_n815), .B2(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n652), .A2(new_n814), .A3(new_n662), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n655), .B1(new_n666), .B2(new_n813), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT110), .B(KEYINPUT55), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n816), .B(new_n256), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n251), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n244), .A2(new_n245), .ZN(new_n826));
  INV_X1    g625(.A(new_n237), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n211), .B1(new_n233), .B2(KEYINPUT17), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n579), .B2(new_n580), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(new_n238), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n826), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT111), .B(new_n827), .C1(new_n829), .C2(new_n238), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n255), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n669), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n807), .B1(new_n824), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n816), .B(new_n836), .C1(new_n822), .C2(new_n823), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n706), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n722), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n670), .A2(new_n257), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n520), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n450), .A2(new_n515), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n675), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n285), .A3(new_n256), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n841), .A2(new_n842), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n450), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT112), .B(new_n686), .C1(new_n841), .C2(new_n842), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n675), .A2(new_n520), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n525), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n256), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n850), .B1(new_n861), .B2(new_n278), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n849), .A2(new_n276), .A3(new_n669), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n669), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G120gat), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(G1341gat));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n564), .A3(new_n691), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n859), .A2(new_n723), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n564), .ZN(G1342gat));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n625), .A3(new_n858), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G134gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n675), .A2(G134gat), .A3(new_n692), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n848), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n876), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n875), .B(new_n878), .C1(new_n846), .C2(new_n847), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  OAI221_X1 g681(.A(new_n874), .B1(new_n875), .B2(new_n877), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT116), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n856), .A2(new_n526), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n686), .A2(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n820), .A2(new_n821), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT117), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n256), .A3(new_n816), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n625), .B1(new_n890), .B2(new_n837), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n577), .B1(new_n891), .B2(new_n840), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n892), .B2(new_n842), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n852), .B2(new_n686), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895), .B2(new_n257), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n450), .A2(new_n518), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n843), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n675), .ZN(new_n899));
  INV_X1    g698(.A(G141gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n256), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g702(.A(G148gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n904), .A3(new_n669), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n839), .A2(new_n692), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n577), .B1(new_n891), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n842), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n686), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n887), .B1(new_n841), .B2(new_n842), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n669), .A3(new_n886), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n895), .A2(new_n744), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(KEYINPUT59), .A3(new_n904), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n905), .B1(new_n915), .B2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n895), .B2(new_n722), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n569), .A3(new_n691), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  NOR4_X1   g720(.A1(new_n898), .A2(G162gat), .A3(new_n675), .A4(new_n692), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT118), .Z(new_n923));
  OAI21_X1  g722(.A(G162gat), .B1(new_n895), .B2(new_n706), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n530), .A2(new_n672), .A3(new_n516), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n853), .B2(new_n854), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n926), .C1(new_n853), .C2(new_n854), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n360), .A3(new_n257), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n845), .A2(new_n675), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT120), .Z(new_n934));
  AOI21_X1  g733(.A(new_n672), .B1(new_n841), .B2(new_n842), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT119), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT121), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n256), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n932), .B1(new_n942), .B2(new_n360), .ZN(G1348gat));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n361), .A3(new_n669), .ZN(new_n944));
  OAI21_X1  g743(.A(G176gat), .B1(new_n931), .B2(new_n744), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  NOR2_X1   g745(.A1(new_n577), .A2(new_n368), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n934), .A2(new_n936), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  OAI21_X1  g748(.A(G183gat), .B1(new_n931), .B2(new_n722), .ZN(new_n950));
  XNOR2_X1  g749(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n949), .A2(new_n956), .A3(new_n950), .A4(new_n951), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(G1350gat));
  NOR2_X1   g757(.A1(new_n706), .A2(G190gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n939), .A2(new_n940), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n928), .A2(new_n625), .A3(new_n930), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(G190gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n961), .B2(G190gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n967), .B(new_n960), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1351gat));
  AND3_X1   g768(.A1(new_n936), .A2(new_n675), .A3(new_n897), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n256), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n675), .A2(new_n526), .A3(new_n520), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT127), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n912), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n256), .A2(G197gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  INV_X1    g775(.A(G204gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n970), .A2(new_n977), .A3(new_n669), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n913), .A2(new_n669), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n970), .A2(new_n342), .A3(new_n691), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n912), .A2(new_n577), .A3(new_n972), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  AOI21_X1  g787(.A(G218gat), .B1(new_n970), .B2(new_n807), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n692), .A2(new_n341), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n989), .B1(new_n974), .B2(new_n990), .ZN(G1355gat));
endmodule


