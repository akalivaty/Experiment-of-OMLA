

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730;

  AND2_X1 U369 ( .A1(n544), .A2(n660), .ZN(n545) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(n500), .Z(n717) );
  INV_X2 U371 ( .A(n631), .ZN(n637) );
  NOR2_X2 U372 ( .A1(n347), .A2(n556), .ZN(n566) );
  NOR2_X2 U373 ( .A1(n554), .A2(KEYINPUT47), .ZN(n347) );
  XNOR2_X2 U374 ( .A(n348), .B(n530), .ZN(n544) );
  NAND2_X2 U375 ( .A1(n418), .A2(n384), .ZN(n348) );
  INV_X2 U376 ( .A(G953), .ZN(n720) );
  NOR2_X1 U377 ( .A1(n660), .A2(n602), .ZN(n626) );
  XOR2_X1 U378 ( .A(G101), .B(G104), .Z(n349) );
  AND2_X1 U379 ( .A1(n363), .A2(n362), .ZN(n609) );
  XNOR2_X1 U380 ( .A(n388), .B(n387), .ZN(n730) );
  BUF_X1 U381 ( .A(n550), .Z(n540) );
  XNOR2_X1 U382 ( .A(n379), .B(n616), .ZN(n415) );
  NAND2_X1 U383 ( .A1(n443), .A2(n441), .ZN(n379) );
  XNOR2_X1 U384 ( .A(n389), .B(n358), .ZN(n681) );
  AND2_X1 U385 ( .A1(n665), .A2(n666), .ZN(n670) );
  XNOR2_X1 U386 ( .A(n403), .B(G143), .ZN(n515) );
  XNOR2_X1 U387 ( .A(G119), .B(G113), .ZN(n448) );
  XNOR2_X2 U388 ( .A(G128), .B(KEYINPUT65), .ZN(n403) );
  XNOR2_X2 U389 ( .A(n419), .B(n498), .ZN(n704) );
  XNOR2_X2 U390 ( .A(n449), .B(n450), .ZN(n419) );
  XOR2_X1 U391 ( .A(G140), .B(G137), .Z(n474) );
  XNOR2_X1 U392 ( .A(n470), .B(G469), .ZN(n546) );
  NOR2_X1 U393 ( .A1(n691), .A2(G902), .ZN(n470) );
  INV_X1 U394 ( .A(KEYINPUT72), .ZN(n530) );
  AND2_X1 U395 ( .A1(n651), .A2(n385), .ZN(n384) );
  XNOR2_X1 U396 ( .A(n428), .B(n516), .ZN(n572) );
  OR2_X1 U397 ( .A1(n699), .A2(G902), .ZN(n428) );
  NOR2_X1 U398 ( .A1(G237), .A2(G953), .ZN(n454) );
  XNOR2_X1 U399 ( .A(n499), .B(n353), .ZN(n468) );
  XOR2_X1 U400 ( .A(KEYINPUT5), .B(G101), .Z(n452) );
  XNOR2_X1 U401 ( .A(G146), .B(G137), .ZN(n451) );
  AND2_X1 U402 ( .A1(n522), .A2(G210), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n446), .B(KEYINPUT74), .ZN(n450) );
  XNOR2_X1 U404 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U405 ( .A(G116), .B(KEYINPUT3), .ZN(n446) );
  XNOR2_X1 U406 ( .A(n474), .B(n468), .ZN(n716) );
  XNOR2_X1 U407 ( .A(n515), .B(n456), .ZN(n499) );
  XNOR2_X1 U408 ( .A(n455), .B(KEYINPUT4), .ZN(n456) );
  INV_X1 U409 ( .A(KEYINPUT64), .ZN(n455) );
  INV_X1 U410 ( .A(n504), .ZN(n463) );
  INV_X1 U411 ( .A(KEYINPUT76), .ZN(n461) );
  NOR2_X1 U412 ( .A1(n580), .A2(n378), .ZN(n395) );
  XNOR2_X1 U413 ( .A(n579), .B(KEYINPUT46), .ZN(n378) );
  INV_X1 U414 ( .A(KEYINPUT44), .ZN(n600) );
  NAND2_X1 U415 ( .A1(n381), .A2(n382), .ZN(n603) );
  INV_X1 U416 ( .A(n654), .ZN(n381) );
  INV_X1 U417 ( .A(KEYINPUT30), .ZN(n434) );
  NOR2_X1 U418 ( .A1(n618), .A2(n411), .ZN(n410) );
  INV_X1 U419 ( .A(G472), .ZN(n411) );
  XNOR2_X1 U420 ( .A(KEYINPUT16), .B(G122), .ZN(n498) );
  XNOR2_X1 U421 ( .A(n400), .B(n397), .ZN(n701) );
  XNOR2_X1 U422 ( .A(n399), .B(n398), .ZN(n397) );
  XNOR2_X1 U423 ( .A(n475), .B(n476), .ZN(n398) );
  XNOR2_X1 U424 ( .A(n425), .B(n424), .ZN(n512) );
  XNOR2_X1 U425 ( .A(G122), .B(KEYINPUT9), .ZN(n424) );
  XNOR2_X1 U426 ( .A(n426), .B(G116), .ZN(n425) );
  XNOR2_X1 U427 ( .A(KEYINPUT103), .B(KEYINPUT7), .ZN(n426) );
  XNOR2_X1 U428 ( .A(n574), .B(n380), .ZN(n680) );
  INV_X1 U429 ( .A(KEYINPUT41), .ZN(n380) );
  XNOR2_X1 U430 ( .A(n433), .B(KEYINPUT39), .ZN(n569) );
  XNOR2_X1 U431 ( .A(n416), .B(n356), .ZN(n598) );
  NOR2_X1 U432 ( .A1(n603), .A2(n365), .ZN(n662) );
  INV_X1 U433 ( .A(KEYINPUT110), .ZN(n548) );
  NAND2_X1 U434 ( .A1(n547), .A2(n382), .ZN(n414) );
  NAND2_X1 U435 ( .A1(n374), .A2(G210), .ZN(n423) );
  INV_X1 U436 ( .A(KEYINPUT73), .ZN(n447) );
  INV_X1 U437 ( .A(KEYINPUT75), .ZN(n460) );
  INV_X1 U438 ( .A(n529), .ZN(n385) );
  OR2_X1 U439 ( .A1(G902), .A2(G237), .ZN(n508) );
  XNOR2_X1 U440 ( .A(G128), .B(KEYINPUT24), .ZN(n476) );
  XNOR2_X1 U441 ( .A(G119), .B(G110), .ZN(n475) );
  XNOR2_X1 U442 ( .A(n477), .B(n474), .ZN(n399) );
  XOR2_X1 U443 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n521) );
  XNOR2_X1 U444 ( .A(G140), .B(G131), .ZN(n520) );
  XNOR2_X1 U445 ( .A(G104), .B(G143), .ZN(n517) );
  XOR2_X1 U446 ( .A(G122), .B(G113), .Z(n518) );
  XNOR2_X1 U447 ( .A(n546), .B(KEYINPUT1), .ZN(n654) );
  INV_X1 U448 ( .A(n651), .ZN(n417) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n487) );
  XNOR2_X1 U450 ( .A(n468), .B(n366), .ZN(n492) );
  XNOR2_X1 U451 ( .A(n453), .B(n368), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U453 ( .A(n463), .B(KEYINPUT93), .ZN(n467) );
  XNOR2_X1 U454 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n581) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n394) );
  NOR2_X1 U457 ( .A1(n608), .A2(n442), .ZN(n441) );
  NOR2_X1 U458 ( .A1(n603), .A2(n614), .ZN(n389) );
  BUF_X1 U459 ( .A(n654), .Z(n396) );
  NAND2_X1 U460 ( .A1(n369), .A2(n639), .ZN(n537) );
  NOR2_X1 U461 ( .A1(n427), .A2(n370), .ZN(n369) );
  OR2_X1 U462 ( .A1(n614), .A2(n551), .ZN(n427) );
  XNOR2_X1 U463 ( .A(n497), .B(KEYINPUT81), .ZN(n542) );
  XNOR2_X1 U464 ( .A(n435), .B(n434), .ZN(n495) );
  NOR2_X1 U465 ( .A1(n550), .A2(n551), .ZN(n553) );
  NAND2_X1 U466 ( .A1(n598), .A2(n396), .ZN(n612) );
  XNOR2_X1 U467 ( .A(n660), .B(KEYINPUT6), .ZN(n614) );
  NAND2_X1 U468 ( .A1(n413), .A2(n410), .ZN(n409) );
  NOR2_X1 U469 ( .A1(n408), .A2(n702), .ZN(n407) );
  NOR2_X1 U470 ( .A1(n413), .A2(n410), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n513), .B(n429), .ZN(n699) );
  XNOR2_X1 U472 ( .A(n515), .B(n514), .ZN(n429) );
  XNOR2_X1 U473 ( .A(G107), .B(G134), .ZN(n511) );
  NOR2_X1 U474 ( .A1(n576), .A2(n680), .ZN(n577) );
  INV_X1 U475 ( .A(KEYINPUT35), .ZN(n401) );
  INV_X1 U476 ( .A(n590), .ZN(n390) );
  INV_X1 U477 ( .A(KEYINPUT32), .ZN(n387) );
  XNOR2_X1 U478 ( .A(n604), .B(n393), .ZN(n642) );
  XNOR2_X1 U479 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n393) );
  XNOR2_X1 U480 ( .A(n570), .B(KEYINPUT108), .ZN(n639) );
  XNOR2_X1 U481 ( .A(n445), .B(KEYINPUT98), .ZN(n602) );
  INV_X1 U482 ( .A(KEYINPUT122), .ZN(n436) );
  NAND2_X1 U483 ( .A1(n431), .A2(n412), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n432), .B(n350), .ZN(n431) );
  INV_X1 U485 ( .A(KEYINPUT56), .ZN(n420) );
  NAND2_X1 U486 ( .A1(n422), .A2(n412), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n423), .B(n359), .ZN(n422) );
  XOR2_X1 U488 ( .A(n697), .B(n361), .Z(n350) );
  INV_X1 U489 ( .A(n653), .ZN(n382) );
  XOR2_X1 U490 ( .A(n494), .B(G472), .Z(n351) );
  AND2_X1 U491 ( .A1(n727), .A2(KEYINPUT70), .ZN(n352) );
  INV_X1 U492 ( .A(n665), .ZN(n551) );
  XNOR2_X1 U493 ( .A(G131), .B(G134), .ZN(n353) );
  AND2_X1 U494 ( .A1(n365), .A2(n418), .ZN(n354) );
  XNOR2_X1 U495 ( .A(n414), .B(KEYINPUT97), .ZN(n601) );
  NOR2_X1 U496 ( .A1(n668), .A2(n417), .ZN(n355) );
  XOR2_X1 U497 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n356) );
  XOR2_X1 U498 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n357) );
  XOR2_X1 U499 ( .A(KEYINPUT89), .B(KEYINPUT33), .Z(n358) );
  XNOR2_X1 U500 ( .A(n690), .B(n689), .ZN(n359) );
  XNOR2_X1 U501 ( .A(KEYINPUT90), .B(n620), .ZN(n702) );
  INV_X1 U502 ( .A(n702), .ZN(n412) );
  XNOR2_X1 U503 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n360) );
  XNOR2_X1 U504 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n361) );
  INV_X1 U505 ( .A(n730), .ZN(n362) );
  NAND2_X1 U506 ( .A1(n592), .A2(n354), .ZN(n363) );
  XNOR2_X1 U507 ( .A(n363), .B(G110), .ZN(G12) );
  NAND2_X1 U508 ( .A1(n375), .A2(n355), .ZN(n416) );
  NAND2_X1 U509 ( .A1(n375), .A2(n601), .ZN(n445) );
  NOR2_X1 U510 ( .A1(n681), .A2(n364), .ZN(n589) );
  INV_X1 U511 ( .A(n375), .ZN(n364) );
  XNOR2_X2 U512 ( .A(n377), .B(n357), .ZN(n375) );
  AND2_X1 U513 ( .A1(n660), .A2(n665), .ZN(n435) );
  INV_X1 U514 ( .A(n660), .ZN(n365) );
  XNOR2_X2 U515 ( .A(n493), .B(n351), .ZN(n660) );
  XNOR2_X1 U516 ( .A(n367), .B(n419), .ZN(n366) );
  NOR2_X1 U517 ( .A1(n537), .A2(n540), .ZN(n538) );
  INV_X1 U518 ( .A(n544), .ZN(n370) );
  NOR2_X2 U519 ( .A1(n648), .A2(n618), .ZN(n374) );
  NAND2_X1 U520 ( .A1(n373), .A2(n371), .ZN(n432) );
  NOR2_X1 U521 ( .A1(n618), .A2(n372), .ZN(n371) );
  INV_X1 U522 ( .A(G475), .ZN(n372) );
  INV_X1 U523 ( .A(n648), .ZN(n373) );
  NAND2_X1 U524 ( .A1(n374), .A2(G217), .ZN(n440) );
  NAND2_X1 U525 ( .A1(n374), .A2(G478), .ZN(n698) );
  NAND2_X1 U526 ( .A1(n374), .A2(G469), .ZN(n694) );
  NAND2_X1 U527 ( .A1(n375), .A2(n662), .ZN(n604) );
  XNOR2_X1 U528 ( .A(n376), .B(n509), .ZN(n550) );
  XNOR2_X1 U529 ( .A(n553), .B(n552), .ZN(n588) );
  NAND2_X1 U530 ( .A1(n688), .A2(n618), .ZN(n376) );
  NAND2_X1 U531 ( .A1(n588), .A2(n587), .ZN(n377) );
  XNOR2_X1 U532 ( .A(n444), .B(n600), .ZN(n443) );
  NAND2_X1 U533 ( .A1(n415), .A2(n719), .ZN(n386) );
  NAND2_X1 U534 ( .A1(n562), .A2(KEYINPUT78), .ZN(n554) );
  AND2_X2 U535 ( .A1(n637), .A2(n606), .ZN(n562) );
  NAND2_X1 U536 ( .A1(n383), .A2(n547), .ZN(n549) );
  XNOR2_X1 U537 ( .A(n545), .B(KEYINPUT28), .ZN(n383) );
  XNOR2_X2 U538 ( .A(n386), .B(n617), .ZN(n648) );
  NAND2_X1 U539 ( .A1(n609), .A2(n352), .ZN(n444) );
  NAND2_X1 U540 ( .A1(n599), .A2(n598), .ZN(n388) );
  NAND2_X1 U541 ( .A1(n391), .A2(n390), .ZN(n402) );
  XNOR2_X1 U542 ( .A(n589), .B(KEYINPUT34), .ZN(n391) );
  NAND2_X1 U543 ( .A1(n392), .A2(n606), .ZN(n607) );
  XNOR2_X1 U544 ( .A(n605), .B(KEYINPUT101), .ZN(n392) );
  XNOR2_X1 U545 ( .A(n479), .B(n717), .ZN(n400) );
  XNOR2_X1 U546 ( .A(n507), .B(n506), .ZN(n688) );
  XNOR2_X1 U547 ( .A(n430), .B(n360), .ZN(G60) );
  XNOR2_X2 U548 ( .A(n402), .B(n401), .ZN(n727) );
  NAND2_X1 U549 ( .A1(n648), .A2(n619), .ZN(n405) );
  NOR2_X1 U550 ( .A1(n406), .A2(n404), .ZN(n622) );
  NAND2_X1 U551 ( .A1(n405), .A2(n407), .ZN(n404) );
  NOR2_X1 U552 ( .A1(n648), .A2(n409), .ZN(n406) );
  INV_X1 U553 ( .A(n619), .ZN(n413) );
  NAND2_X1 U554 ( .A1(n496), .A2(n601), .ZN(n497) );
  NAND2_X1 U555 ( .A1(n593), .A2(n651), .ZN(n653) );
  NAND2_X1 U556 ( .A1(n415), .A2(n720), .ZN(n712) );
  NAND2_X1 U557 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U558 ( .A(n593), .ZN(n418) );
  NOR2_X2 U559 ( .A1(G902), .A2(n701), .ZN(n484) );
  XNOR2_X1 U560 ( .A(n421), .B(n420), .ZN(G51) );
  NAND2_X1 U561 ( .A1(n569), .A2(n570), .ZN(n571) );
  NAND2_X1 U562 ( .A1(n542), .A2(n666), .ZN(n433) );
  XNOR2_X1 U563 ( .A(n437), .B(n436), .ZN(G66) );
  NAND2_X1 U564 ( .A1(n438), .A2(n412), .ZN(n437) );
  XNOR2_X1 U565 ( .A(n440), .B(n439), .ZN(n438) );
  INV_X1 U566 ( .A(n701), .ZN(n439) );
  NAND2_X1 U567 ( .A1(n611), .A2(n623), .ZN(n442) );
  INV_X1 U568 ( .A(KEYINPUT85), .ZN(n557) );
  XNOR2_X1 U569 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U570 ( .A(n501), .B(KEYINPUT18), .ZN(n502) );
  INV_X1 U571 ( .A(KEYINPUT71), .ZN(n567) );
  XNOR2_X1 U572 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U573 ( .A(n505), .B(n463), .ZN(n506) );
  INV_X1 U574 ( .A(n396), .ZN(n595) );
  INV_X1 U575 ( .A(KEYINPUT63), .ZN(n621) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n458) );
  XNOR2_X1 U577 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U578 ( .A(n454), .B(KEYINPUT80), .ZN(n522) );
  XNOR2_X1 U579 ( .A(n492), .B(KEYINPUT113), .ZN(n457) );
  XNOR2_X1 U580 ( .A(n458), .B(n457), .ZN(n619) );
  XNOR2_X1 U581 ( .A(G110), .B(G107), .ZN(n459) );
  XNOR2_X1 U582 ( .A(n349), .B(n459), .ZN(n703) );
  XNOR2_X1 U583 ( .A(n703), .B(n462), .ZN(n504) );
  NAND2_X1 U584 ( .A1(G227), .A2(n720), .ZN(n465) );
  XNOR2_X1 U585 ( .A(G146), .B(KEYINPUT82), .ZN(n464) );
  XNOR2_X1 U586 ( .A(n469), .B(n716), .ZN(n691) );
  XOR2_X1 U587 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n473) );
  XNOR2_X2 U588 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  NAND2_X1 U589 ( .A1(G234), .A2(n618), .ZN(n471) );
  XNOR2_X1 U590 ( .A(KEYINPUT20), .B(n471), .ZN(n480) );
  NAND2_X1 U591 ( .A1(n480), .A2(G221), .ZN(n472) );
  XNOR2_X1 U592 ( .A(n473), .B(n472), .ZN(n651) );
  XOR2_X2 U593 ( .A(G125), .B(G146), .Z(n500) );
  XOR2_X1 U594 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n477) );
  NAND2_X1 U595 ( .A1(G234), .A2(n720), .ZN(n478) );
  XOR2_X1 U596 ( .A(KEYINPUT8), .B(n478), .Z(n510) );
  NAND2_X1 U597 ( .A1(G221), .A2(n510), .ZN(n479) );
  XOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n482) );
  NAND2_X1 U599 ( .A1(n480), .A2(G217), .ZN(n481) );
  XNOR2_X1 U600 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X2 U601 ( .A(n484), .B(n483), .ZN(n593) );
  NOR2_X1 U602 ( .A1(G900), .A2(n720), .ZN(n485) );
  NAND2_X1 U603 ( .A1(G902), .A2(n485), .ZN(n486) );
  NAND2_X1 U604 ( .A1(G952), .A2(n720), .ZN(n583) );
  NAND2_X1 U605 ( .A1(n486), .A2(n583), .ZN(n490) );
  XOR2_X1 U606 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n488) );
  XNOR2_X1 U607 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U608 ( .A(KEYINPUT79), .B(n489), .Z(n585) );
  INV_X1 U609 ( .A(n585), .ZN(n649) );
  NAND2_X1 U610 ( .A1(n490), .A2(n649), .ZN(n529) );
  NAND2_X1 U611 ( .A1(n508), .A2(G214), .ZN(n491) );
  XOR2_X1 U612 ( .A(n491), .B(KEYINPUT91), .Z(n665) );
  XNOR2_X1 U613 ( .A(KEYINPUT77), .B(KEYINPUT99), .ZN(n494) );
  NOR2_X1 U614 ( .A1(G902), .A2(n492), .ZN(n493) );
  NOR2_X1 U615 ( .A1(n529), .A2(n495), .ZN(n496) );
  XNOR2_X1 U616 ( .A(n704), .B(n499), .ZN(n507) );
  XOR2_X1 U617 ( .A(n500), .B(KEYINPUT17), .Z(n503) );
  NAND2_X1 U618 ( .A1(G224), .A2(n720), .ZN(n501) );
  NAND2_X1 U619 ( .A1(G210), .A2(n508), .ZN(n509) );
  XNOR2_X1 U620 ( .A(KEYINPUT38), .B(n540), .ZN(n666) );
  NAND2_X1 U621 ( .A1(n510), .A2(G217), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U623 ( .A(KEYINPUT104), .B(G478), .ZN(n516) );
  INV_X1 U624 ( .A(n572), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U626 ( .A(n717), .B(n519), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n521), .B(n520), .ZN(n524) );
  NAND2_X1 U628 ( .A1(n522), .A2(G214), .ZN(n523) );
  XOR2_X1 U629 ( .A(n524), .B(n523), .Z(n525) );
  XNOR2_X1 U630 ( .A(n526), .B(n525), .ZN(n697) );
  NOR2_X1 U631 ( .A1(G902), .A2(n697), .ZN(n528) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(G475), .ZN(n527) );
  XNOR2_X1 U633 ( .A(n528), .B(n527), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT102), .ZN(n532) );
  NOR2_X1 U635 ( .A1(n533), .A2(n532), .ZN(n641) );
  NAND2_X1 U636 ( .A1(n569), .A2(n641), .ZN(n646) );
  NAND2_X1 U637 ( .A1(n533), .A2(n532), .ZN(n543) );
  INV_X1 U638 ( .A(n543), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT109), .B(n537), .ZN(n534) );
  NAND2_X1 U640 ( .A1(n534), .A2(n396), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n535), .B(KEYINPUT43), .ZN(n536) );
  NAND2_X1 U642 ( .A1(n536), .A2(n540), .ZN(n647) );
  NAND2_X1 U643 ( .A1(n646), .A2(n647), .ZN(n582) );
  XNOR2_X1 U644 ( .A(KEYINPUT36), .B(n538), .ZN(n539) );
  NAND2_X1 U645 ( .A1(n539), .A2(n595), .ZN(n645) );
  NAND2_X1 U646 ( .A1(n573), .A2(n572), .ZN(n590) );
  NOR2_X1 U647 ( .A1(n540), .A2(n590), .ZN(n541) );
  NAND2_X1 U648 ( .A1(n542), .A2(n541), .ZN(n636) );
  NAND2_X1 U649 ( .A1(n645), .A2(n636), .ZN(n556) );
  INV_X1 U650 ( .A(n641), .ZN(n630) );
  NAND2_X1 U651 ( .A1(n630), .A2(n543), .ZN(n669) );
  XNOR2_X1 U652 ( .A(KEYINPUT86), .B(n669), .ZN(n606) );
  INV_X1 U653 ( .A(n546), .ZN(n547) );
  XNOR2_X2 U654 ( .A(n549), .B(n548), .ZN(n575) );
  XOR2_X1 U655 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n552) );
  NAND2_X1 U656 ( .A1(n575), .A2(n588), .ZN(n631) );
  NAND2_X1 U657 ( .A1(n631), .A2(KEYINPUT47), .ZN(n558) );
  XNOR2_X1 U658 ( .A(n558), .B(n557), .ZN(n561) );
  NAND2_X1 U659 ( .A1(KEYINPUT78), .A2(n669), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n559), .A2(KEYINPUT47), .ZN(n560) );
  NAND2_X1 U661 ( .A1(n561), .A2(n560), .ZN(n564) );
  NOR2_X1 U662 ( .A1(n562), .A2(KEYINPUT78), .ZN(n563) );
  NOR2_X1 U663 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U664 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U665 ( .A(n568), .B(n567), .ZN(n580) );
  XNOR2_X2 U666 ( .A(n571), .B(KEYINPUT40), .ZN(n729) );
  XNOR2_X1 U667 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n578) );
  NOR2_X1 U668 ( .A1(n573), .A2(n572), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n670), .A2(n591), .ZN(n574) );
  INV_X1 U670 ( .A(n575), .ZN(n576) );
  XNOR2_X1 U671 ( .A(n578), .B(n577), .ZN(n728) );
  NAND2_X1 U672 ( .A1(n729), .A2(n728), .ZN(n579) );
  NOR2_X2 U673 ( .A1(n582), .A2(n581), .ZN(n719) );
  NOR2_X1 U674 ( .A1(G898), .A2(n720), .ZN(n706) );
  NAND2_X1 U675 ( .A1(G902), .A2(n706), .ZN(n584) );
  AND2_X1 U676 ( .A1(n584), .A2(n583), .ZN(n586) );
  NOR2_X1 U677 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U678 ( .A(n591), .ZN(n668) );
  XNOR2_X1 U679 ( .A(n612), .B(KEYINPUT107), .ZN(n592) );
  XOR2_X1 U680 ( .A(n593), .B(KEYINPUT106), .Z(n613) );
  INV_X1 U681 ( .A(n613), .ZN(n650) );
  XOR2_X1 U682 ( .A(KEYINPUT84), .B(n614), .Z(n594) );
  NOR2_X1 U683 ( .A1(n650), .A2(n594), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U685 ( .A(KEYINPUT83), .B(n597), .ZN(n599) );
  NOR2_X1 U686 ( .A1(n626), .A2(n642), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT105), .ZN(n608) );
  NOR2_X1 U688 ( .A1(KEYINPUT70), .A2(n727), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n623) );
  XOR2_X1 U691 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n616) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n617) );
  NOR2_X1 U693 ( .A1(G952), .A2(n720), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(G57) );
  XNOR2_X1 U695 ( .A(G101), .B(KEYINPUT114), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(G3) );
  NAND2_X1 U697 ( .A1(n639), .A2(n626), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U700 ( .A1(n626), .A2(n641), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(G107), .B(n629), .ZN(G9) );
  NOR2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n633) );
  XNOR2_X1 U705 ( .A(G128), .B(KEYINPUT116), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(G30) );
  XNOR2_X1 U708 ( .A(G143), .B(n636), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n639), .A2(n637), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(G146), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n642), .A2(n639), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(G113), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(G116), .ZN(G18) );
  XOR2_X1 U715 ( .A(G125), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(G27) );
  XNOR2_X1 U717 ( .A(G134), .B(n646), .ZN(G36) );
  XNOR2_X1 U718 ( .A(G140), .B(n647), .ZN(G42) );
  NAND2_X1 U719 ( .A1(n720), .A2(n648), .ZN(n686) );
  NAND2_X1 U720 ( .A1(G952), .A2(n649), .ZN(n679) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(KEYINPUT49), .B(n652), .ZN(n658) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n656) );
  NAND2_X1 U724 ( .A1(n396), .A2(n653), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U729 ( .A(KEYINPUT51), .B(n663), .Z(n664) );
  NOR2_X1 U730 ( .A1(n680), .A2(n664), .ZN(n676) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U734 ( .A(KEYINPUT118), .B(n671), .Z(n672) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n674), .A2(n681), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U738 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n684), .B(KEYINPUT119), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U744 ( .A(KEYINPUT53), .B(n687), .ZN(G75) );
  XOR2_X1 U745 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n690) );
  XNOR2_X1 U746 ( .A(n688), .B(KEYINPUT55), .ZN(n689) );
  XNOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U751 ( .A1(n702), .A2(n696), .ZN(G54) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n702), .A2(n700), .ZN(G63) );
  XOR2_X1 U754 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U755 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U756 ( .A(KEYINPUT125), .B(n707), .Z(n715) );
  XOR2_X1 U757 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n709) );
  NAND2_X1 U758 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U760 ( .A1(G898), .A2(n710), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n711), .B(KEYINPUT124), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U764 ( .A(n716), .B(n717), .Z(n718) );
  XOR2_X1 U765 ( .A(KEYINPUT126), .B(n718), .Z(n722) );
  XOR2_X1 U766 ( .A(n722), .B(n719), .Z(n721) );
  NAND2_X1 U767 ( .A1(n721), .A2(n720), .ZN(n726) );
  XNOR2_X1 U768 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U769 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U770 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U772 ( .A(n727), .B(G122), .ZN(G24) );
  XNOR2_X1 U773 ( .A(G137), .B(n728), .ZN(G39) );
  XNOR2_X1 U774 ( .A(n729), .B(G131), .ZN(G33) );
  XOR2_X1 U775 ( .A(G119), .B(n730), .Z(G21) );
endmodule

