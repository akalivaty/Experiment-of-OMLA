

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n432, n433, n434, n435, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804;

  XNOR2_X1 U371 ( .A(n619), .B(KEYINPUT38), .ZN(n749) );
  NOR2_X2 U372 ( .A1(n647), .A2(n420), .ZN(n563) );
  AND2_X2 U373 ( .A1(n768), .A2(n754), .ZN(n615) );
  NAND2_X2 U374 ( .A1(n350), .A2(n569), .ZN(n571) );
  NOR2_X2 U375 ( .A1(n568), .A2(n761), .ZN(n350) );
  XNOR2_X2 U376 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X2 U377 ( .A1(n351), .A2(n435), .ZN(n601) );
  AND2_X2 U378 ( .A1(n437), .A2(n439), .ZN(n351) );
  NAND2_X1 U379 ( .A1(n632), .A2(n631), .ZN(n353) );
  XNOR2_X2 U380 ( .A(n394), .B(KEYINPUT40), .ZN(n632) );
  XNOR2_X2 U381 ( .A(n352), .B(KEYINPUT82), .ZN(n605) );
  NAND2_X2 U382 ( .A1(n599), .A2(n598), .ZN(n352) );
  XOR2_X2 U383 ( .A(n484), .B(n483), .Z(n485) );
  AND2_X2 U384 ( .A1(n417), .A2(n416), .ZN(n415) );
  XNOR2_X2 U385 ( .A(n353), .B(n633), .ZN(n393) );
  NOR2_X2 U386 ( .A1(n645), .A2(n624), .ZN(n625) );
  XNOR2_X2 U387 ( .A(n549), .B(n541), .ZN(n686) );
  XNOR2_X2 U388 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X2 U389 ( .A1(n415), .A2(n420), .ZN(n384) );
  XNOR2_X2 U390 ( .A(n549), .B(n548), .ZN(n711) );
  AND2_X2 U391 ( .A1(n461), .A2(n463), .ZN(n460) );
  AND2_X2 U392 ( .A1(n403), .A2(n577), .ZN(n583) );
  OR2_X2 U393 ( .A1(n686), .A2(G902), .ZN(n542) );
  NAND2_X2 U394 ( .A1(n354), .A2(n387), .ZN(n665) );
  AND2_X2 U395 ( .A1(n389), .A2(n388), .ZN(n354) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n535) );
  XNOR2_X1 U397 ( .A(G113), .B(G143), .ZN(n521) );
  AND2_X2 U398 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X2 U399 ( .A1(n368), .A2(n466), .ZN(n464) );
  NOR2_X2 U400 ( .A1(n777), .A2(n735), .ZN(n630) );
  XNOR2_X2 U401 ( .A(n564), .B(n543), .ZN(n568) );
  XNOR2_X2 U402 ( .A(n542), .B(G472), .ZN(n564) );
  NOR2_X1 U403 ( .A1(n572), .A2(n773), .ZN(n588) );
  INV_X1 U404 ( .A(n720), .ZN(n447) );
  AND2_X1 U405 ( .A1(n444), .A2(n442), .ZN(n432) );
  AND2_X1 U406 ( .A1(n443), .A2(n573), .ZN(n442) );
  NOR2_X1 U407 ( .A1(n584), .A2(n429), .ZN(n428) );
  INV_X1 U408 ( .A(KEYINPUT0), .ZN(n356) );
  NOR2_X1 U409 ( .A1(n788), .A2(n667), .ZN(n738) );
  AND2_X1 U410 ( .A1(n391), .A2(n660), .ZN(n388) );
  NOR2_X1 U411 ( .A1(n705), .A2(n596), .ZN(n597) );
  NAND2_X1 U412 ( .A1(n432), .A2(n357), .ZN(n435) );
  XNOR2_X1 U413 ( .A(n428), .B(KEYINPUT32), .ZN(n707) );
  NOR2_X1 U414 ( .A1(n584), .A2(n471), .ZN(n585) );
  NOR2_X1 U415 ( .A1(n757), .A2(n399), .ZN(n621) );
  XNOR2_X1 U416 ( .A(n513), .B(n512), .ZN(n592) );
  XNOR2_X1 U417 ( .A(G140), .B(KEYINPUT10), .ZN(n422) );
  INV_X1 U418 ( .A(G953), .ZN(n499) );
  XNOR2_X2 U419 ( .A(n498), .B(n356), .ZN(n355) );
  INV_X2 U420 ( .A(n355), .ZN(n572) );
  XNOR2_X1 U421 ( .A(n486), .B(n485), .ZN(n618) );
  XNOR2_X2 U422 ( .A(n449), .B(n453), .ZN(n794) );
  XNOR2_X2 U423 ( .A(n508), .B(n454), .ZN(n453) );
  XNOR2_X2 U424 ( .A(n540), .B(n546), .ZN(n449) );
  AND2_X2 U425 ( .A1(n425), .A2(n430), .ZN(n708) );
  NOR2_X1 U426 ( .A1(n603), .A2(KEYINPUT44), .ZN(n604) );
  INV_X1 U427 ( .A(KEYINPUT111), .ZN(n379) );
  XNOR2_X1 U428 ( .A(n500), .B(KEYINPUT8), .ZN(n554) );
  NAND2_X1 U429 ( .A1(n390), .A2(n392), .ZN(n387) );
  INV_X1 U430 ( .A(n738), .ZN(n430) );
  XNOR2_X1 U431 ( .A(n562), .B(n358), .ZN(n421) );
  AND2_X1 U432 ( .A1(n709), .A2(n414), .ZN(n418) );
  INV_X1 U433 ( .A(G134), .ZN(n504) );
  NAND2_X1 U434 ( .A1(n604), .A2(n469), .ZN(n467) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n491) );
  NAND2_X1 U436 ( .A1(G469), .A2(n414), .ZN(n413) );
  NAND2_X1 U437 ( .A1(n550), .A2(G902), .ZN(n416) );
  XNOR2_X1 U438 ( .A(G116), .B(KEYINPUT98), .ZN(n537) );
  OR2_X1 U439 ( .A1(n554), .A2(n501), .ZN(n503) );
  INV_X1 U440 ( .A(KEYINPUT77), .ZN(n445) );
  XNOR2_X1 U441 ( .A(G101), .B(G107), .ZN(n545) );
  NOR2_X1 U442 ( .A1(n652), .A2(n655), .ZN(n402) );
  INV_X1 U443 ( .A(KEYINPUT36), .ZN(n401) );
  OR2_X1 U444 ( .A1(n448), .A2(n569), .ZN(n471) );
  XNOR2_X1 U445 ( .A(n560), .B(n559), .ZN(n709) );
  NOR2_X1 U446 ( .A1(n457), .A2(n606), .ZN(n456) );
  INV_X1 U447 ( .A(n467), .ZN(n457) );
  INV_X1 U448 ( .A(KEYINPUT109), .ZN(n408) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  NAND2_X1 U450 ( .A1(n434), .A2(n433), .ZN(n444) );
  NOR2_X1 U451 ( .A1(n572), .A2(KEYINPUT34), .ZN(n433) );
  INV_X1 U452 ( .A(G237), .ZN(n482) );
  XNOR2_X1 U453 ( .A(n424), .B(n423), .ZN(n561) );
  NAND2_X1 U454 ( .A1(n606), .A2(G234), .ZN(n423) );
  XNOR2_X1 U455 ( .A(n528), .B(KEYINPUT95), .ZN(n424) );
  XOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT20), .Z(n528) );
  XOR2_X1 U457 ( .A(G122), .B(G104), .Z(n522) );
  XOR2_X1 U458 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n515) );
  XOR2_X1 U459 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n517) );
  NAND2_X1 U460 ( .A1(n380), .A2(n378), .ZN(n377) );
  XNOR2_X1 U461 ( .A(n627), .B(KEYINPUT1), .ZN(n567) );
  INV_X1 U462 ( .A(KEYINPUT16), .ZN(n454) );
  XNOR2_X1 U463 ( .A(G128), .B(G137), .ZN(n555) );
  XNOR2_X1 U464 ( .A(G110), .B(G119), .ZN(n556) );
  XNOR2_X1 U465 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n552) );
  XNOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n551) );
  NAND2_X1 U467 ( .A1(n362), .A2(n455), .ZN(n788) );
  INV_X1 U468 ( .A(KEYINPUT79), .ZN(n661) );
  XNOR2_X1 U469 ( .A(n494), .B(KEYINPUT91), .ZN(n782) );
  XNOR2_X1 U470 ( .A(n506), .B(n400), .ZN(n668) );
  XNOR2_X1 U471 ( .A(n534), .B(n510), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n397), .B(n544), .ZN(n547) );
  XNOR2_X1 U473 ( .A(n545), .B(G140), .ZN(n397) );
  XNOR2_X1 U474 ( .A(n371), .B(n370), .ZN(n800) );
  INV_X1 U475 ( .A(KEYINPUT113), .ZN(n370) );
  NOR2_X1 U476 ( .A1(n646), .A2(n647), .ZN(n371) );
  BUF_X1 U477 ( .A(n601), .Z(n706) );
  INV_X1 U478 ( .A(KEYINPUT81), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n710) );
  INV_X1 U480 ( .A(n709), .ZN(n409) );
  NAND2_X1 U481 ( .A1(n367), .A2(G217), .ZN(n410) );
  INV_X1 U482 ( .A(KEYINPUT56), .ZN(n404) );
  AND2_X1 U483 ( .A1(n441), .A2(KEYINPUT35), .ZN(n357) );
  INV_X1 U484 ( .A(n420), .ZN(n766) );
  BUF_X1 U485 ( .A(n499), .Z(n677) );
  XOR2_X1 U486 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n358) );
  INV_X1 U487 ( .A(n765), .ZN(n419) );
  INV_X1 U488 ( .A(n754), .ZN(n399) );
  XOR2_X1 U489 ( .A(n490), .B(KEYINPUT19), .Z(n359) );
  AND2_X1 U490 ( .A1(n751), .A2(n419), .ZN(n360) );
  BUF_X2 U491 ( .A(n567), .Z(n762) );
  AND2_X1 U492 ( .A1(n468), .A2(n456), .ZN(n361) );
  AND2_X1 U493 ( .A1(n468), .A2(n467), .ZN(n362) );
  INV_X1 U494 ( .A(G902), .ZN(n414) );
  XOR2_X1 U495 ( .A(n366), .B(n693), .Z(n363) );
  XNOR2_X1 U496 ( .A(KEYINPUT124), .B(n668), .ZN(n364) );
  NAND2_X1 U497 ( .A1(n664), .A2(KEYINPUT2), .ZN(n365) );
  INV_X1 U498 ( .A(KEYINPUT78), .ZN(n470) );
  NOR2_X1 U499 ( .A1(n677), .A2(G952), .ZN(n717) );
  NAND2_X1 U500 ( .A1(n375), .A2(n447), .ZN(n394) );
  NAND2_X1 U501 ( .A1(n468), .A2(n456), .ZN(n465) );
  BUF_X1 U502 ( .A(n619), .Z(n655) );
  BUF_X2 U503 ( .A(n564), .Z(n768) );
  XNOR2_X1 U504 ( .A(n762), .B(KEYINPUT84), .ZN(n647) );
  XNOR2_X1 U505 ( .A(n740), .B(KEYINPUT69), .ZN(n662) );
  INV_X1 U506 ( .A(n568), .ZN(n448) );
  AND2_X1 U507 ( .A1(n447), .A2(n398), .ZN(n446) );
  BUF_X1 U508 ( .A(n694), .Z(n366) );
  NAND2_X1 U509 ( .A1(n605), .A2(n469), .ZN(n468) );
  AND2_X2 U510 ( .A1(n425), .A2(n430), .ZN(n367) );
  XNOR2_X1 U511 ( .A(n632), .B(G131), .ZN(G33) );
  BUF_X1 U512 ( .A(n464), .Z(n455) );
  AND2_X1 U513 ( .A1(n464), .A2(KEYINPUT78), .ZN(n459) );
  INV_X1 U514 ( .A(n605), .ZN(n368) );
  NOR2_X1 U515 ( .A1(n645), .A2(n399), .ZN(n398) );
  XNOR2_X2 U516 ( .A(n418), .B(n421), .ZN(n420) );
  AND2_X2 U517 ( .A1(n601), .A2(KEYINPUT64), .ZN(n575) );
  INV_X1 U518 ( .A(n464), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n372), .B(n359), .ZN(n635) );
  NOR2_X2 U520 ( .A1(n618), .A2(n399), .ZN(n372) );
  NOR2_X1 U521 ( .A1(n373), .A2(n719), .ZN(n595) );
  NAND2_X1 U522 ( .A1(n373), .A2(n728), .ZN(n673) );
  NAND2_X1 U523 ( .A1(n373), .A2(n447), .ZN(n674) );
  XNOR2_X1 U524 ( .A(n588), .B(n374), .ZN(n373) );
  INV_X1 U525 ( .A(KEYINPUT31), .ZN(n374) );
  NAND2_X1 U526 ( .A1(n375), .A2(n728), .ZN(n672) );
  XNOR2_X2 U527 ( .A(n620), .B(KEYINPUT39), .ZN(n375) );
  NAND2_X1 U528 ( .A1(n376), .A2(KEYINPUT111), .ZN(n382) );
  INV_X1 U529 ( .A(n411), .ZN(n376) );
  NAND2_X1 U530 ( .A1(n380), .A2(n411), .ZN(n607) );
  NAND2_X1 U531 ( .A1(n381), .A2(n377), .ZN(n385) );
  AND2_X1 U532 ( .A1(n411), .A2(n379), .ZN(n378) );
  INV_X1 U533 ( .A(n384), .ZN(n380) );
  NAND2_X1 U534 ( .A1(n384), .A2(KEYINPUT111), .ZN(n383) );
  NAND2_X1 U535 ( .A1(n385), .A2(n622), .ZN(n614) );
  NAND2_X1 U536 ( .A1(n393), .A2(n386), .ZN(n389) );
  AND2_X1 U537 ( .A1(n649), .A2(n651), .ZN(n386) );
  INV_X1 U538 ( .A(n393), .ZN(n390) );
  OR2_X1 U539 ( .A1(n649), .A2(n651), .ZN(n391) );
  INV_X1 U540 ( .A(n651), .ZN(n392) );
  INV_X1 U541 ( .A(n554), .ZN(n407) );
  NAND2_X1 U542 ( .A1(n462), .A2(n470), .ZN(n461) );
  AND2_X2 U543 ( .A1(n395), .A2(n420), .ZN(n705) );
  XNOR2_X1 U544 ( .A(n585), .B(n396), .ZN(n395) );
  AND2_X2 U545 ( .A1(n412), .A2(n419), .ZN(n411) );
  NAND2_X1 U546 ( .A1(n361), .A2(n459), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n402), .B(n401), .ZN(n646) );
  NAND2_X1 U548 ( .A1(n575), .A2(n602), .ZN(n403) );
  XNOR2_X1 U549 ( .A(n405), .B(n404), .ZN(G51) );
  NAND2_X1 U550 ( .A1(n696), .A2(n670), .ZN(n405) );
  XNOR2_X1 U551 ( .A(n406), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U552 ( .A1(n671), .A2(n670), .ZN(n406) );
  NAND2_X1 U553 ( .A1(n407), .A2(G221), .ZN(n558) );
  XNOR2_X1 U554 ( .A(n794), .B(n481), .ZN(n694) );
  XNOR2_X1 U555 ( .A(n597), .B(n408), .ZN(n598) );
  NAND2_X1 U556 ( .A1(n420), .A2(n419), .ZN(n761) );
  NAND2_X1 U557 ( .A1(n415), .A2(n412), .ZN(n627) );
  OR2_X2 U558 ( .A1(n711), .A2(n413), .ZN(n412) );
  NAND2_X1 U559 ( .A1(n711), .A2(n550), .ZN(n417) );
  XNOR2_X2 U560 ( .A(n520), .B(n422), .ZN(n676) );
  XNOR2_X2 U561 ( .A(G146), .B(G125), .ZN(n520) );
  NAND2_X1 U562 ( .A1(n426), .A2(n365), .ZN(n425) );
  XNOR2_X1 U563 ( .A(n427), .B(n445), .ZN(n426) );
  NAND2_X1 U564 ( .A1(n663), .A2(n662), .ZN(n427) );
  NAND2_X1 U565 ( .A1(n563), .A2(n568), .ZN(n429) );
  XNOR2_X2 U566 ( .A(n530), .B(KEYINPUT22), .ZN(n584) );
  INV_X1 U567 ( .A(n760), .ZN(n434) );
  NAND2_X1 U568 ( .A1(n438), .A2(n574), .ZN(n437) );
  NAND2_X1 U569 ( .A1(n442), .A2(n441), .ZN(n438) );
  NAND2_X1 U570 ( .A1(n440), .A2(n574), .ZN(n439) );
  INV_X1 U571 ( .A(n444), .ZN(n440) );
  NAND2_X1 U572 ( .A1(n760), .A2(KEYINPUT34), .ZN(n441) );
  NAND2_X1 U573 ( .A1(n572), .A2(KEYINPUT34), .ZN(n443) );
  NAND2_X1 U574 ( .A1(n448), .A2(n446), .ZN(n652) );
  NAND2_X1 U575 ( .A1(n465), .A2(n470), .ZN(n463) );
  XNOR2_X2 U576 ( .A(n450), .B(G110), .ZN(n546) );
  XNOR2_X2 U577 ( .A(G104), .B(KEYINPUT87), .ZN(n450) );
  XNOR2_X2 U578 ( .A(n452), .B(n451), .ZN(n540) );
  XNOR2_X2 U579 ( .A(G119), .B(KEYINPUT3), .ZN(n451) );
  XNOR2_X2 U580 ( .A(G101), .B(G113), .ZN(n452) );
  XNOR2_X2 U581 ( .A(n472), .B(G107), .ZN(n508) );
  NAND2_X1 U582 ( .A1(n460), .A2(n458), .ZN(n663) );
  NOR2_X1 U583 ( .A1(n604), .A2(n469), .ZN(n466) );
  INV_X1 U584 ( .A(KEYINPUT45), .ZN(n469) );
  XNOR2_X2 U585 ( .A(G116), .B(G122), .ZN(n472) );
  INV_X1 U586 ( .A(n803), .ZN(n631) );
  INV_X1 U587 ( .A(n717), .ZN(n670) );
  XNOR2_X2 U588 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n520), .B(n532), .ZN(n476) );
  XNOR2_X1 U590 ( .A(KEYINPUT72), .B(KEYINPUT17), .ZN(n474) );
  XNOR2_X1 U591 ( .A(KEYINPUT18), .B(KEYINPUT71), .ZN(n473) );
  XNOR2_X1 U592 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n476), .B(n475), .ZN(n480) );
  NAND2_X1 U594 ( .A1(n499), .A2(G224), .ZN(n477) );
  XNOR2_X1 U595 ( .A(n477), .B(KEYINPUT88), .ZN(n478) );
  XNOR2_X2 U596 ( .A(G143), .B(G128), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n505), .B(n478), .ZN(n479) );
  XNOR2_X1 U598 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U599 ( .A(n606), .ZN(n664) );
  NOR2_X1 U600 ( .A1(n694), .A2(n664), .ZN(n486) );
  NAND2_X1 U601 ( .A1(n414), .A2(n482), .ZN(n487) );
  NAND2_X1 U602 ( .A1(n487), .A2(G210), .ZN(n484) );
  INV_X1 U603 ( .A(KEYINPUT73), .ZN(n483) );
  NAND2_X1 U604 ( .A1(n487), .A2(G214), .ZN(n489) );
  INV_X1 U605 ( .A(KEYINPUT89), .ZN(n488) );
  XNOR2_X1 U606 ( .A(n489), .B(n488), .ZN(n754) );
  INV_X1 U607 ( .A(KEYINPUT65), .ZN(n490) );
  XOR2_X1 U608 ( .A(KEYINPUT90), .B(KEYINPUT14), .Z(n492) );
  XNOR2_X1 U609 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U610 ( .A(KEYINPUT68), .B(n493), .Z(n495) );
  NAND2_X1 U611 ( .A1(n495), .A2(G952), .ZN(n494) );
  NAND2_X1 U612 ( .A1(n782), .A2(n677), .ZN(n611) );
  NAND2_X1 U613 ( .A1(G902), .A2(n495), .ZN(n608) );
  XOR2_X1 U614 ( .A(G898), .B(KEYINPUT92), .Z(n791) );
  NAND2_X1 U615 ( .A1(G953), .A2(n791), .ZN(n795) );
  OR2_X1 U616 ( .A1(n608), .A2(n795), .ZN(n496) );
  NAND2_X1 U617 ( .A1(n611), .A2(n496), .ZN(n497) );
  NAND2_X1 U618 ( .A1(n635), .A2(n497), .ZN(n498) );
  NAND2_X1 U619 ( .A1(n499), .A2(G234), .ZN(n500) );
  INV_X1 U620 ( .A(G217), .ZN(n501) );
  XOR2_X1 U621 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U622 ( .A(n503), .B(n502), .ZN(n506) );
  XNOR2_X2 U623 ( .A(n505), .B(n504), .ZN(n534) );
  XNOR2_X1 U624 ( .A(KEYINPUT104), .B(KEYINPUT7), .ZN(n507) );
  XNOR2_X1 U625 ( .A(n507), .B(KEYINPUT9), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n508), .B(n509), .ZN(n510) );
  NAND2_X1 U627 ( .A1(n668), .A2(n414), .ZN(n513) );
  XNOR2_X1 U628 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U629 ( .A(n511), .B(G478), .ZN(n512) );
  NAND2_X1 U630 ( .A1(G214), .A2(n535), .ZN(n514) );
  XNOR2_X1 U631 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U632 ( .A(G131), .B(KEYINPUT12), .ZN(n516) );
  XNOR2_X1 U633 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U634 ( .A(n519), .B(n518), .Z(n525) );
  XNOR2_X1 U635 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U636 ( .A(n676), .B(n523), .ZN(n524) );
  XNOR2_X1 U637 ( .A(n525), .B(n524), .ZN(n699) );
  NAND2_X1 U638 ( .A1(n699), .A2(n414), .ZN(n527) );
  XNOR2_X1 U639 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  XNOR2_X1 U640 ( .A(n527), .B(n526), .ZN(n591) );
  AND2_X1 U641 ( .A1(n592), .A2(n591), .ZN(n751) );
  NAND2_X1 U642 ( .A1(n561), .A2(G221), .ZN(n529) );
  XNOR2_X1 U643 ( .A(n529), .B(KEYINPUT21), .ZN(n765) );
  NAND2_X1 U644 ( .A1(n355), .A2(n360), .ZN(n530) );
  XNOR2_X1 U645 ( .A(G131), .B(G137), .ZN(n531) );
  XNOR2_X1 U646 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X2 U647 ( .A(n534), .B(n533), .ZN(n675) );
  XNOR2_X2 U648 ( .A(n675), .B(G146), .ZN(n549) );
  NAND2_X1 U649 ( .A1(n535), .A2(G210), .ZN(n536) );
  XNOR2_X1 U650 ( .A(n536), .B(KEYINPUT5), .ZN(n538) );
  XNOR2_X1 U651 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U652 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U653 ( .A(KEYINPUT108), .B(KEYINPUT6), .ZN(n543) );
  NAND2_X1 U654 ( .A1(n677), .A2(G227), .ZN(n544) );
  XNOR2_X1 U655 ( .A(n547), .B(n546), .ZN(n548) );
  INV_X1 U656 ( .A(G469), .ZN(n550) );
  XNOR2_X1 U657 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U658 ( .A(n676), .B(n553), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U660 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U661 ( .A1(n561), .A2(G217), .ZN(n562) );
  NOR2_X1 U662 ( .A1(n768), .A2(n420), .ZN(n565) );
  NAND2_X1 U663 ( .A1(n762), .A2(n565), .ZN(n566) );
  NOR2_X1 U664 ( .A1(n584), .A2(n566), .ZN(n684) );
  NOR2_X2 U665 ( .A1(n707), .A2(n684), .ZN(n602) );
  INV_X1 U666 ( .A(n567), .ZN(n569) );
  INV_X1 U667 ( .A(KEYINPUT33), .ZN(n570) );
  XNOR2_X2 U668 ( .A(n571), .B(n570), .ZN(n760) );
  OR2_X1 U669 ( .A1(n591), .A2(n592), .ZN(n640) );
  INV_X1 U670 ( .A(n640), .ZN(n573) );
  INV_X1 U671 ( .A(KEYINPUT35), .ZN(n574) );
  INV_X1 U672 ( .A(KEYINPUT64), .ZN(n576) );
  OR2_X1 U673 ( .A1(n576), .A2(KEYINPUT44), .ZN(n577) );
  INV_X1 U674 ( .A(n602), .ZN(n581) );
  INV_X1 U675 ( .A(n601), .ZN(n579) );
  NAND2_X1 U676 ( .A1(n576), .A2(KEYINPUT44), .ZN(n578) );
  NOR2_X1 U677 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U678 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U679 ( .A1(n583), .A2(n582), .ZN(n599) );
  INV_X1 U680 ( .A(n761), .ZN(n586) );
  NAND2_X1 U681 ( .A1(n768), .A2(n586), .ZN(n587) );
  OR2_X1 U682 ( .A1(n762), .A2(n587), .ZN(n773) );
  OR2_X1 U683 ( .A1(n607), .A2(n768), .ZN(n589) );
  NOR2_X1 U684 ( .A1(n572), .A2(n589), .ZN(n719) );
  INV_X1 U685 ( .A(n592), .ZN(n590) );
  NAND2_X1 U686 ( .A1(n590), .A2(n591), .ZN(n723) );
  INV_X1 U687 ( .A(n591), .ZN(n593) );
  NAND2_X1 U688 ( .A1(n593), .A2(n592), .ZN(n720) );
  NAND2_X1 U689 ( .A1(n723), .A2(n720), .ZN(n594) );
  XNOR2_X1 U690 ( .A(n594), .B(KEYINPUT107), .ZN(n748) );
  NOR2_X1 U691 ( .A1(n595), .A2(n748), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n602), .A2(n706), .ZN(n603) );
  NOR2_X1 U693 ( .A1(G900), .A2(n608), .ZN(n609) );
  NAND2_X1 U694 ( .A1(G953), .A2(n609), .ZN(n610) );
  NAND2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U696 ( .A(n612), .B(KEYINPUT74), .ZN(n622) );
  INV_X1 U697 ( .A(KEYINPUT70), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n614), .B(n613), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n615), .B(KEYINPUT30), .ZN(n616) );
  AND2_X2 U700 ( .A1(n617), .A2(n616), .ZN(n642) );
  BUF_X1 U701 ( .A(n618), .Z(n619) );
  NAND2_X1 U702 ( .A1(n642), .A2(n749), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n749), .A2(n751), .ZN(n757) );
  XNOR2_X1 U704 ( .A(n621), .B(KEYINPUT41), .ZN(n777) );
  AND2_X1 U705 ( .A1(n622), .A2(n419), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n623), .A2(n766), .ZN(n645) );
  INV_X1 U707 ( .A(n768), .ZN(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(KEYINPUT28), .ZN(n629) );
  INV_X1 U709 ( .A(KEYINPUT112), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n735) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT42), .ZN(n803) );
  INV_X1 U713 ( .A(KEYINPUT46), .ZN(n633) );
  BUF_X1 U714 ( .A(n635), .Z(n636) );
  INV_X1 U715 ( .A(n636), .ZN(n637) );
  OR2_X1 U716 ( .A1(n748), .A2(n637), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n735), .A2(n638), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n639), .B(KEYINPUT47), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n655), .A2(n640), .ZN(n641) );
  AND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n733) );
  INV_X1 U721 ( .A(n733), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n648), .A2(n800), .ZN(n649) );
  INV_X1 U724 ( .A(KEYINPUT80), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT48), .ZN(n651) );
  INV_X1 U726 ( .A(n723), .ZN(n728) );
  INV_X1 U727 ( .A(n652), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n762), .A2(n653), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT43), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n658) );
  INV_X1 U731 ( .A(KEYINPUT110), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n804) );
  INV_X1 U733 ( .A(n804), .ZN(n659) );
  AND2_X1 U734 ( .A1(n672), .A2(n659), .ZN(n660) );
  XNOR2_X2 U735 ( .A(n665), .B(n661), .ZN(n740) );
  INV_X1 U736 ( .A(n665), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n367), .A2(G478), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(n364), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(G134), .ZN(G36) );
  XNOR2_X1 U741 ( .A(n673), .B(G116), .ZN(G18) );
  XNOR2_X1 U742 ( .A(n674), .B(G113), .ZN(G15) );
  XOR2_X1 U743 ( .A(n675), .B(n676), .Z(n679) );
  XNOR2_X1 U744 ( .A(n740), .B(n679), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n683) );
  XNOR2_X1 U746 ( .A(n679), .B(G227), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n680), .A2(G900), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n681), .A2(G953), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(G72) );
  XOR2_X1 U750 ( .A(G110), .B(n684), .Z(G12) );
  NAND2_X1 U751 ( .A1(n708), .A2(G472), .ZN(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X2 U754 ( .A1(n689), .A2(n717), .ZN(n691) );
  XOR2_X1 U755 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n690) );
  XNOR2_X1 U756 ( .A(n691), .B(n690), .ZN(G57) );
  NAND2_X1 U757 ( .A1(n367), .A2(G210), .ZN(n695) );
  XNOR2_X1 U758 ( .A(KEYINPUT83), .B(KEYINPUT54), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT55), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n695), .B(n363), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n708), .A2(G475), .ZN(n701) );
  XNOR2_X1 U762 ( .A(KEYINPUT85), .B(KEYINPUT123), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT59), .ZN(n698) );
  XNOR2_X1 U764 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X2 U765 ( .A1(n702), .A2(n717), .ZN(n704) );
  XNOR2_X1 U766 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n703) );
  XNOR2_X1 U767 ( .A(n704), .B(n703), .ZN(G60) );
  XOR2_X1 U768 ( .A(n705), .B(G101), .Z(G3) );
  XNOR2_X1 U769 ( .A(n706), .B(G122), .ZN(G24) );
  XOR2_X1 U770 ( .A(n707), .B(G119), .Z(G21) );
  NOR2_X1 U771 ( .A1(n710), .A2(n717), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n367), .A2(G469), .ZN(n716) );
  XOR2_X1 U773 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n713) );
  XNOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n712) );
  XOR2_X1 U775 ( .A(n713), .B(n712), .Z(n714) );
  XNOR2_X1 U776 ( .A(n711), .B(n714), .ZN(n715) );
  XNOR2_X1 U777 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(G54) );
  INV_X1 U779 ( .A(n719), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n724), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(G104), .B(KEYINPUT115), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(G6) );
  NOR2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n725) );
  XNOR2_X1 U785 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U786 ( .A(G107), .B(n727), .ZN(G9) );
  NAND2_X1 U787 ( .A1(n636), .A2(n728), .ZN(n729) );
  NOR2_X1 U788 ( .A1(n735), .A2(n729), .ZN(n731) );
  XNOR2_X1 U789 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n730) );
  XNOR2_X1 U790 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U791 ( .A(G128), .B(n732), .ZN(G30) );
  XOR2_X1 U792 ( .A(G143), .B(n733), .Z(G45) );
  NAND2_X1 U793 ( .A1(n636), .A2(n447), .ZN(n734) );
  NOR2_X1 U794 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U795 ( .A(G146), .B(n736), .Z(G48) );
  XNOR2_X1 U796 ( .A(KEYINPUT2), .B(KEYINPUT75), .ZN(n743) );
  AND2_X1 U797 ( .A1(n740), .A2(n743), .ZN(n737) );
  NOR2_X1 U798 ( .A1(n737), .A2(KEYINPUT76), .ZN(n739) );
  NOR2_X1 U799 ( .A1(n739), .A2(n738), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n740), .A2(KEYINPUT76), .ZN(n742) );
  INV_X1 U801 ( .A(n788), .ZN(n741) );
  NAND2_X1 U802 ( .A1(n742), .A2(n741), .ZN(n744) );
  NAND2_X1 U803 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U804 ( .A1(n746), .A2(n745), .ZN(n786) );
  NOR2_X1 U805 ( .A1(n777), .A2(n760), .ZN(n747) );
  NOR2_X1 U806 ( .A1(G953), .A2(n747), .ZN(n784) );
  INV_X1 U807 ( .A(n748), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n750), .A2(n749), .ZN(n753) );
  INV_X1 U809 ( .A(n751), .ZN(n752) );
  NAND2_X1 U810 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U811 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U812 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U813 ( .A(KEYINPUT120), .B(n758), .Z(n759) );
  NOR2_X1 U814 ( .A1(n760), .A2(n759), .ZN(n779) );
  NAND2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(KEYINPUT119), .ZN(n764) );
  XNOR2_X1 U817 ( .A(n764), .B(KEYINPUT50), .ZN(n772) );
  NAND2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n767), .B(KEYINPUT49), .ZN(n769) );
  OR2_X1 U820 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n770), .B(KEYINPUT118), .ZN(n771) );
  OR2_X1 U822 ( .A1(n772), .A2(n771), .ZN(n774) );
  AND2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U824 ( .A(KEYINPUT51), .B(n775), .Z(n776) );
  NOR2_X1 U825 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U826 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U827 ( .A(KEYINPUT52), .B(n780), .Z(n781) );
  NAND2_X1 U828 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U829 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U830 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U831 ( .A(KEYINPUT53), .B(n787), .ZN(G75) );
  NOR2_X1 U832 ( .A1(n788), .A2(G953), .ZN(n793) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n789) );
  XOR2_X1 U834 ( .A(KEYINPUT61), .B(n789), .Z(n790) );
  NOR2_X1 U835 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U836 ( .A1(n793), .A2(n792), .ZN(n799) );
  XOR2_X1 U837 ( .A(KEYINPUT126), .B(n794), .Z(n796) );
  NAND2_X1 U838 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U839 ( .A(n797), .B(KEYINPUT127), .ZN(n798) );
  XOR2_X1 U840 ( .A(n799), .B(n798), .Z(G69) );
  XOR2_X1 U841 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n802) );
  XNOR2_X1 U842 ( .A(n800), .B(G125), .ZN(n801) );
  XNOR2_X1 U843 ( .A(n802), .B(n801), .ZN(G27) );
  XOR2_X1 U844 ( .A(n803), .B(G137), .Z(G39) );
  XOR2_X1 U845 ( .A(G140), .B(n804), .Z(G42) );
endmodule

