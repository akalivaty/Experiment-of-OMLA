//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n207), .B2(KEYINPUT83), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n209), .A3(new_n206), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n208), .A2(new_n210), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218));
  INV_X1    g017(.A(new_n206), .ZN(new_n219));
  NOR2_X1   g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT83), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n210), .A3(KEYINPUT15), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT84), .A2(KEYINPUT15), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT84), .A2(KEYINPUT15), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n214), .A2(new_n216), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n217), .A2(new_n218), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n218), .A3(new_n222), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT17), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n218), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n222), .A2(new_n234), .A3(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n229), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G8gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G15gat), .B(G22gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(G1gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n243), .B2(KEYINPUT86), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(G1gat), .B2(new_n241), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT87), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n248), .B1(new_n228), .B2(new_n230), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n253), .A4(new_n254), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n228), .A2(new_n230), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n252), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n258), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G141gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G197gat), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT11), .B(G169gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n271), .A3(new_n258), .A4(new_n265), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(KEYINPUT22), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G211gat), .B(G218gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(G155gat), .B2(G162gat), .ZN(new_n287));
  INV_X1    g086(.A(G155gat), .ZN(new_n288));
  INV_X1    g087(.A(G162gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI22_X1  g089(.A1(new_n285), .A2(new_n287), .B1(KEYINPUT76), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G155gat), .B(G162gat), .Z(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n284), .A2(new_n296), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n293), .B1(new_n298), .B2(new_n294), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G78gat), .B(G106gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(G22gat), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT31), .B(G50gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n292), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n291), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(KEYINPUT1), .B2(new_n314), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n312), .A2(new_n313), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n321), .A2(new_n323), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT4), .B1(new_n293), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n291), .A2(new_n292), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n291), .A2(new_n292), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT3), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n295), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n293), .A2(new_n326), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n324), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT39), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT79), .B(KEYINPUT39), .C1(new_n339), .C2(new_n335), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT0), .ZN(new_n346));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g147(.A(KEYINPUT39), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n349), .A3(new_n335), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT40), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n348), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n328), .A2(new_n355), .A3(new_n334), .A4(new_n332), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n313), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n293), .A2(new_n326), .A3(KEYINPUT4), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n332), .A2(new_n358), .A3(new_n334), .A4(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n339), .B2(new_n335), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n356), .A2(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n357), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n354), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n344), .A2(KEYINPUT40), .A3(new_n348), .A4(new_n350), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n353), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT27), .B(G183gat), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n369), .A2(KEYINPUT68), .ZN(new_n370));
  INV_X1    g169(.A(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(KEYINPUT68), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(KEYINPUT28), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT28), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n378), .A2(KEYINPUT26), .ZN(new_n379));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n378), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  OR2_X1    g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n378), .A2(KEYINPUT23), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(G169gat), .B2(G176gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n380), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n387), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT64), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT64), .B(new_n387), .C1(new_n392), .C2(new_n396), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n396), .A2(new_n387), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n388), .A2(KEYINPUT66), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n388), .A2(KEYINPUT66), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n389), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n391), .B(KEYINPUT65), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n368), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n368), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(KEYINPUT29), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n284), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND3_X1  g219(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(new_n284), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n386), .A2(new_n413), .A3(new_n407), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n420), .A4(new_n424), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n420), .B(KEYINPUT75), .ZN(new_n429));
  INV_X1    g228(.A(new_n424), .ZN(new_n430));
  INV_X1    g229(.A(new_n411), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n410), .B1(new_n386), .B2(new_n407), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n413), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n422), .B1(new_n433), .B2(new_n415), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n427), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n310), .B1(new_n367), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n417), .A2(new_n439), .A3(new_n424), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT37), .B1(new_n430), .B2(new_n434), .ZN(new_n441));
  INV_X1    g240(.A(new_n420), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n443), .B2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n429), .A2(new_n438), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n421), .A2(new_n284), .A3(new_n423), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n284), .B1(new_n433), .B2(new_n415), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT80), .B1(new_n452), .B2(new_n440), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n417), .A2(new_n439), .A3(new_n424), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n422), .B1(new_n412), .B2(new_n416), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(KEYINPUT37), .A3(new_n449), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n448), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n357), .B1(new_n360), .B2(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n360), .A2(new_n361), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n348), .A3(new_n363), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n365), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT6), .B(new_n354), .C1(new_n362), .C2(new_n364), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n465), .A2(new_n466), .A3(new_n425), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n437), .B1(new_n447), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n386), .A2(new_n407), .A3(new_n326), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n326), .B1(new_n386), .B2(new_n407), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT32), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G71gat), .B(G99gat), .Z(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(KEYINPUT32), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n470), .B2(KEYINPUT72), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n472), .A2(new_n473), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n470), .ZN(new_n493));
  NOR4_X1   g292(.A1(new_n472), .A2(new_n473), .A3(new_n471), .A4(new_n490), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n495), .B(new_n481), .C1(new_n486), .C2(new_n487), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n486), .A2(new_n487), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(KEYINPUT73), .A3(new_n495), .A4(new_n481), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(KEYINPUT36), .A3(new_n499), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n465), .A2(new_n466), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n436), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n427), .A2(new_n428), .A3(new_n435), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n465), .A2(new_n466), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n310), .A3(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n469), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT35), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n503), .B2(new_n500), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n309), .A3(new_n499), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n508), .A2(new_n507), .A3(new_n436), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT78), .B1(new_n510), .B2(new_n511), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n522), .B2(KEYINPUT35), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n277), .B1(new_n514), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n509), .B2(new_n512), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n500), .A2(new_n503), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n469), .A2(new_n506), .A3(new_n513), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT82), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n276), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT41), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n533), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G99gat), .B(G106gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT8), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(G85gat), .B(G92gat), .C1(KEYINPUT91), .C2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g351(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n541), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n542), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n560));
  AND2_X1   g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n559), .A2(new_n562), .A3(new_n540), .A4(new_n547), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n565), .B(new_n541), .C1(new_n551), .C2(new_n555), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n571), .A2(new_n259), .B1(new_n535), .B2(new_n534), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n571), .A2(new_n574), .B1(new_n231), .B2(new_n238), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(KEYINPUT94), .A3(new_n570), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT95), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n566), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT93), .B1(new_n564), .B2(new_n566), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n239), .A2(new_n580), .A3(new_n576), .A4(KEYINPUT95), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n539), .B(new_n573), .C1(new_n577), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT96), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n239), .A2(new_n580), .A3(new_n576), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n572), .B1(new_n587), .B2(new_n581), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n539), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(KEYINPUT97), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n573), .B1(new_n577), .B2(new_n582), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n538), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT97), .B1(new_n584), .B2(new_n590), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n537), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n584), .A2(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(KEYINPUT98), .A3(new_n538), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n588), .B2(new_n539), .ZN(new_n601));
  INV_X1    g400(.A(new_n537), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT9), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT89), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  OR2_X1    g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G57gat), .A2(G64gat), .ZN(new_n610));
  OR2_X1    g409(.A1(G57gat), .A2(G64gat), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n611), .B(new_n610), .C1(new_n605), .C2(KEYINPUT9), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n608), .A3(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT20), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n619), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n249), .B1(new_n616), .B2(new_n615), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n596), .A2(new_n604), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n596), .A2(new_n604), .A3(new_n631), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n556), .A2(new_n563), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT100), .B1(new_n634), .B2(new_n615), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n564), .A2(new_n566), .A3(new_n615), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n613), .B(new_n609), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n556), .A4(new_n563), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT101), .Z(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n615), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n569), .A2(new_n570), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n635), .A2(new_n636), .A3(new_n639), .A4(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n641), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n644), .A2(new_n654), .A3(new_n650), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n532), .A2(KEYINPUT102), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT82), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT82), .B1(new_n529), .B2(new_n530), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n275), .B(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n508), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND4_X1  g468(.A1(new_n666), .A2(KEYINPUT42), .A3(new_n436), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n666), .A2(new_n436), .A3(new_n669), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n240), .B1(new_n666), .B2(new_n436), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n672), .B1(new_n673), .B2(new_n677), .ZN(G1325gat));
  NOR2_X1   g477(.A1(new_n528), .A2(G15gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n666), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n506), .B1(new_n660), .B2(new_n665), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1326gat));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n666), .B2(new_n310), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n666), .A2(new_n687), .A3(new_n310), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT105), .B(new_n309), .C1(new_n660), .C2(new_n665), .ZN(new_n692));
  INV_X1    g491(.A(new_n686), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n694), .ZN(G1327gat));
  XOR2_X1   g494(.A(new_n658), .B(KEYINPUT106), .Z(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n276), .A3(new_n628), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n596), .A2(new_n604), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n661), .B2(new_n662), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n529), .B2(new_n530), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT107), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n699), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n698), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n511), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n598), .A2(new_n603), .ZN(new_n711));
  INV_X1    g510(.A(new_n595), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n591), .A3(new_n593), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n713), .B2(new_n537), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n628), .A3(new_n658), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n532), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n508), .A2(new_n215), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n716), .A2(new_n710), .A3(new_n717), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n718), .A3(new_n719), .ZN(G1328gat));
  OAI21_X1  g519(.A(G36gat), .B1(new_n708), .B2(new_n510), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n436), .A2(new_n211), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT46), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  OR3_X1    g522(.A1(new_n716), .A2(KEYINPUT46), .A3(new_n722), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AND4_X1   g525(.A1(new_n203), .A2(new_n532), .A3(new_n527), .A4(new_n715), .ZN(new_n727));
  INV_X1    g526(.A(new_n506), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n524), .A2(new_n531), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n704), .B1(new_n729), .B2(new_n699), .ZN(new_n730));
  INV_X1    g529(.A(new_n705), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n699), .A2(new_n704), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n702), .A3(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n728), .B(new_n697), .C1(new_n730), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n727), .B1(new_n734), .B2(G43gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n726), .B1(new_n735), .B2(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n203), .B1(new_n707), .B2(new_n728), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n737), .B(KEYINPUT47), .C1(new_n738), .C2(new_n727), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n736), .A2(new_n739), .ZN(G1330gat));
  NOR3_X1   g539(.A1(new_n716), .A2(G50gat), .A3(new_n309), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n310), .B(new_n697), .C1(new_n730), .C2(new_n733), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n204), .B1(new_n707), .B2(new_n310), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n742), .B1(new_n749), .B2(new_n741), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1331gat));
  NOR2_X1   g550(.A1(new_n731), .A2(new_n702), .ZN(new_n752));
  INV_X1    g551(.A(new_n696), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n633), .A2(new_n275), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n511), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT110), .B(G57gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  OAI22_X1  g557(.A1(new_n755), .A2(new_n510), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT49), .B(G64gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n752), .A2(new_n436), .A3(new_n754), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT111), .Z(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n755), .B2(new_n506), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n528), .A2(G71gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n755), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g566(.A1(new_n755), .A2(new_n309), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT112), .B(G78gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n628), .A2(new_n275), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n658), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n701), .B2(new_n706), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n511), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n699), .B(new_n771), .C1(new_n514), .C2(new_n523), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT51), .ZN(new_n777));
  INV_X1    g576(.A(new_n658), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n508), .A2(new_n548), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NOR2_X1   g580(.A1(new_n777), .A2(new_n753), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n549), .A3(new_n436), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n549), .B1(new_n773), .B2(new_n436), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n785), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(new_n783), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n774), .B2(new_n506), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n528), .A2(G99gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n779), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g592(.A(G106gat), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n773), .B2(new_n310), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n309), .A2(G106gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n796), .A2(KEYINPUT113), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n801), .B2(new_n795), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n630), .A2(new_n276), .A3(new_n632), .A4(new_n778), .ZN(new_n804));
  INV_X1    g603(.A(new_n628), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n647), .A2(new_n642), .A3(new_n648), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT114), .A4(new_n642), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n650), .A3(KEYINPUT54), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n654), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n657), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n657), .A3(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n810), .A2(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n817), .A2(new_n275), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n253), .B1(new_n250), .B2(new_n254), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n823), .A2(KEYINPUT116), .B1(new_n261), .B2(new_n264), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n270), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n658), .A2(new_n826), .A3(new_n274), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(new_n596), .A3(new_n604), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n826), .A2(new_n274), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n818), .A3(new_n817), .A4(new_n821), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n596), .B2(new_n604), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n805), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n310), .B1(new_n804), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n511), .A2(new_n436), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n527), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n276), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n511), .B1(new_n804), .B2(new_n833), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n519), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n436), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n275), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n837), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n836), .A2(new_n319), .A3(new_n753), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n658), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n319), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n841), .A2(new_n847), .A3(new_n628), .ZN(new_n848));
  OAI21_X1  g647(.A(G127gat), .B1(new_n836), .B2(new_n805), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  OR4_X1    g649(.A1(G134gat), .A2(new_n840), .A3(new_n436), .A4(new_n714), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n836), .B2(new_n714), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n506), .A2(new_n835), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n309), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n810), .A2(new_n860), .A3(new_n813), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n820), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n815), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(KEYINPUT118), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n275), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT118), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n827), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n714), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n699), .A2(new_n830), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n628), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n804), .B1(new_n871), .B2(KEYINPUT119), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(new_n628), .C1(new_n868), .C2(new_n870), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n858), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n804), .A2(new_n833), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n310), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n857), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n276), .B(new_n856), .C1(new_n875), .C2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(G141gat), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n728), .A2(new_n309), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n839), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n883), .A2(new_n880), .A3(new_n275), .A4(new_n510), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n879), .B2(new_n880), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI221_X1 g686(.A(new_n884), .B1(KEYINPUT120), .B2(KEYINPUT58), .C1(new_n879), .C2(new_n880), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(G1344gat));
  AND2_X1   g688(.A1(new_n883), .A2(new_n510), .ZN(new_n890));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n658), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n858), .ZN(new_n894));
  INV_X1    g693(.A(new_n871), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n309), .B1(new_n895), .B2(new_n804), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n778), .B1(new_n856), .B2(KEYINPUT121), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n897), .B(new_n898), .C1(KEYINPUT121), .C2(new_n856), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n856), .B1(new_n875), .B2(new_n878), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n891), .C1(new_n901), .C2(new_n658), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n890), .A2(new_n288), .A3(new_n628), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n901), .A2(new_n628), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n288), .ZN(G1346gat));
  NAND4_X1  g705(.A1(new_n883), .A2(new_n289), .A3(new_n510), .A4(new_n699), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n901), .A2(new_n699), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n289), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n508), .A2(new_n510), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n876), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n519), .ZN(new_n912));
  AOI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n275), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n527), .A2(new_n910), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT122), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n834), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n834), .A2(KEYINPUT123), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n275), .A2(G169gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n920), .B2(new_n753), .ZN(new_n924));
  INV_X1    g723(.A(G176gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n912), .A2(new_n925), .A3(new_n658), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1349gat));
  OAI21_X1  g726(.A(G183gat), .B1(new_n920), .B2(new_n805), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n628), .A2(new_n370), .A3(new_n372), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n932), .B(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n912), .A2(new_n371), .A3(new_n699), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n699), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(G190gat), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n937), .B2(G190gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  AND2_X1   g740(.A1(new_n506), .A2(new_n910), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n897), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(new_n944), .A3(new_n276), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n911), .A2(new_n882), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n275), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n949), .A3(new_n658), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n943), .B2(new_n753), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n946), .A2(new_n279), .A3(new_n628), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n897), .A2(new_n628), .A3(new_n942), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n943), .B2(new_n714), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n946), .A2(new_n280), .A3(new_n699), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


