

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G2104), .A2(n514), .ZN(n857) );
  NOR2_X2 U550 ( .A1(n586), .A2(n585), .ZN(G164) );
  NOR2_X2 U551 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  OR2_X1 U552 ( .A1(n611), .A2(n593), .ZN(n595) );
  NOR2_X1 U553 ( .A1(n924), .A2(n632), .ZN(n634) );
  NAND2_X1 U554 ( .A1(n689), .A2(n691), .ZN(n611) );
  NOR2_X1 U555 ( .A1(n662), .A2(n661), .ZN(n678) );
  AND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n689) );
  INV_X1 U557 ( .A(KEYINPUT83), .ZN(n583) );
  INV_X1 U558 ( .A(KEYINPUT27), .ZN(n594) );
  XNOR2_X1 U559 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n633) );
  NOR2_X1 U561 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U562 ( .A(KEYINPUT32), .ZN(n675) );
  XNOR2_X1 U563 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U564 ( .A1(G651), .A2(n555), .ZN(n790) );
  AND2_X1 U565 ( .A1(n514), .A2(G2104), .ZN(n862) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n786) );
  INV_X1 U567 ( .A(G2105), .ZN(n514) );
  NAND2_X1 U568 ( .A1(n862), .A2(G101), .ZN(n513) );
  XOR2_X1 U569 ( .A(KEYINPUT23), .B(n513), .Z(n516) );
  NAND2_X1 U570 ( .A1(n857), .A2(G125), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U572 ( .A(n517), .B(KEYINPUT64), .ZN(n523) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n518), .Z(n865) );
  NAND2_X1 U574 ( .A1(G137), .A2(n865), .ZN(n520) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n858) );
  NAND2_X1 U576 ( .A1(G113), .A2(n858), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U578 ( .A(KEYINPUT65), .B(n521), .Z(n522) );
  NOR2_X2 U579 ( .A1(n523), .A2(n522), .ZN(G160) );
  INV_X1 U580 ( .A(G651), .ZN(n527) );
  NOR2_X1 U581 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n524), .Z(n785) );
  NAND2_X1 U583 ( .A1(G64), .A2(n785), .ZN(n526) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n555) );
  NAND2_X1 U585 ( .A1(G52), .A2(n790), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n555), .A2(n527), .ZN(n789) );
  NAND2_X1 U588 ( .A1(G77), .A2(n789), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G90), .A2(n786), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n530), .Z(n531) );
  NOR2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U593 ( .A(KEYINPUT67), .B(n533), .Z(G171) );
  INV_X1 U594 ( .A(G171), .ZN(G301) );
  NAND2_X1 U595 ( .A1(G63), .A2(n785), .ZN(n535) );
  NAND2_X1 U596 ( .A1(G51), .A2(n790), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U598 ( .A(KEYINPUT6), .B(n536), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n786), .A2(G89), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT4), .ZN(n539) );
  NAND2_X1 U601 ( .A1(G76), .A2(n789), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT5), .B(n540), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT73), .B(n541), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G75), .A2(n789), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G88), .A2(n786), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G62), .A2(n785), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G50), .A2(n790), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(G166) );
  NAND2_X1 U615 ( .A1(G49), .A2(n790), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G74), .A2(G651), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT76), .B(n553), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n785), .A2(n554), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n555), .A2(G87), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(G288) );
  INV_X1 U622 ( .A(G166), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G61), .A2(n785), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G86), .A2(n786), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT77), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G48), .A2(n790), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n789), .A2(G73), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT2), .B(n563), .Z(n564) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT78), .B(n566), .Z(G305) );
  NAND2_X1 U633 ( .A1(G60), .A2(n785), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G47), .A2(n790), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G72), .A2(n789), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT66), .B(n569), .Z(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n786), .A2(G85), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(G290) );
  NAND2_X1 U641 ( .A1(G138), .A2(n865), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G102), .A2(n862), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n574) );
  NAND2_X1 U644 ( .A1(KEYINPUT84), .A2(n574), .ZN(n580) );
  INV_X1 U645 ( .A(KEYINPUT84), .ZN(n578) );
  AND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G126), .A2(n857), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G114), .A2(n858), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n691) );
  BUF_X2 U654 ( .A(n611), .Z(n666) );
  NAND2_X1 U655 ( .A1(G8), .A2(n666), .ZN(n730) );
  NOR2_X1 U656 ( .A1(G1966), .A2(n730), .ZN(n662) );
  NAND2_X1 U657 ( .A1(G65), .A2(n785), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G53), .A2(n790), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G78), .A2(n789), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G91), .A2(n786), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n924) );
  INV_X1 U664 ( .A(KEYINPUT90), .ZN(n599) );
  INV_X1 U665 ( .A(G2072), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G1956), .A2(n666), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n599), .B(n598), .ZN(n632) );
  NAND2_X1 U669 ( .A1(n924), .A2(n632), .ZN(n631) );
  NAND2_X1 U670 ( .A1(n785), .A2(G56), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT14), .ZN(n607) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(KEYINPUT70), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n786), .A2(G81), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT12), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G68), .A2(n789), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT71), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G43), .A2(n790), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n936) );
  INV_X1 U682 ( .A(n611), .ZN(n639) );
  AND2_X1 U683 ( .A1(n639), .A2(G1996), .ZN(n612) );
  XOR2_X1 U684 ( .A(n612), .B(KEYINPUT26), .Z(n614) );
  NAND2_X1 U685 ( .A1(n666), .A2(G1341), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U687 ( .A1(n936), .A2(n615), .ZN(n626) );
  NAND2_X1 U688 ( .A1(G79), .A2(n789), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G54), .A2(n790), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G66), .A2(n785), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G92), .A2(n786), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT15), .ZN(n921) );
  NAND2_X1 U696 ( .A1(G1348), .A2(n666), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G2067), .A2(n639), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n921), .A2(n627), .ZN(n625) );
  OR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n921), .A2(n627), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT29), .ZN(n643) );
  XNOR2_X1 U707 ( .A(G2078), .B(KEYINPUT89), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(KEYINPUT25), .ZN(n952) );
  NOR2_X1 U709 ( .A1(n952), .A2(n666), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n639), .A2(G1961), .ZN(n640) );
  NOR2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n647) );
  NOR2_X1 U712 ( .A1(G301), .A2(n647), .ZN(n642) );
  NOR2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n652) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n666), .ZN(n658) );
  NOR2_X1 U715 ( .A1(n662), .A2(n658), .ZN(n644) );
  NAND2_X1 U716 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U717 ( .A(KEYINPUT30), .B(n645), .ZN(n646) );
  NOR2_X1 U718 ( .A1(G168), .A2(n646), .ZN(n649) );
  AND2_X1 U719 ( .A1(G301), .A2(n647), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT31), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT91), .ZN(n664) );
  INV_X1 U723 ( .A(n664), .ZN(n655) );
  INV_X1 U724 ( .A(KEYINPUT92), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n664), .A2(KEYINPUT92), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n658), .A2(G8), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U730 ( .A1(G286), .A2(G8), .ZN(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n674) );
  INV_X1 U732 ( .A(G8), .ZN(n672) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n730), .ZN(n665) );
  XNOR2_X1 U734 ( .A(KEYINPUT93), .B(n665), .ZN(n669) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n666), .ZN(n667) );
  NOR2_X1 U736 ( .A1(G166), .A2(n667), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT94), .ZN(n671) );
  OR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  AND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n721) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n928) );
  INV_X1 U743 ( .A(n928), .ZN(n681) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(KEYINPUT95), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n721), .A2(n682), .ZN(n685) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n929) );
  INV_X1 U749 ( .A(n929), .ZN(n683) );
  OR2_X1 U750 ( .A1(n683), .A2(n730), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n686), .A2(KEYINPUT33), .ZN(n720) );
  NAND2_X1 U753 ( .A1(n928), .A2(KEYINPUT33), .ZN(n687) );
  OR2_X1 U754 ( .A1(n687), .A2(n730), .ZN(n688) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n939) );
  NAND2_X1 U756 ( .A1(n688), .A2(n939), .ZN(n718) );
  INV_X1 U757 ( .A(n689), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n753) );
  XNOR2_X1 U759 ( .A(KEYINPUT37), .B(G2067), .ZN(n741) );
  NAND2_X1 U760 ( .A1(G104), .A2(n862), .ZN(n693) );
  NAND2_X1 U761 ( .A1(G140), .A2(n865), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U763 ( .A(KEYINPUT34), .B(n694), .ZN(n699) );
  NAND2_X1 U764 ( .A1(G128), .A2(n857), .ZN(n696) );
  NAND2_X1 U765 ( .A1(G116), .A2(n858), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT35), .B(n697), .Z(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U769 ( .A(KEYINPUT36), .B(n700), .ZN(n873) );
  NOR2_X1 U770 ( .A1(n741), .A2(n873), .ZN(n984) );
  NAND2_X1 U771 ( .A1(n753), .A2(n984), .ZN(n751) );
  NAND2_X1 U772 ( .A1(G105), .A2(n862), .ZN(n701) );
  XNOR2_X1 U773 ( .A(n701), .B(KEYINPUT38), .ZN(n708) );
  NAND2_X1 U774 ( .A1(G129), .A2(n857), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G141), .A2(n865), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U777 ( .A1(n858), .A2(G117), .ZN(n704) );
  XOR2_X1 U778 ( .A(KEYINPUT86), .B(n704), .Z(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n844) );
  AND2_X1 U781 ( .A1(n844), .A2(G1996), .ZN(n974) );
  NAND2_X1 U782 ( .A1(n865), .A2(G131), .ZN(n711) );
  NAND2_X1 U783 ( .A1(G95), .A2(n862), .ZN(n709) );
  XOR2_X1 U784 ( .A(KEYINPUT85), .B(n709), .Z(n710) );
  NAND2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U786 ( .A1(G119), .A2(n857), .ZN(n713) );
  NAND2_X1 U787 ( .A1(G107), .A2(n858), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n872) );
  AND2_X1 U790 ( .A1(n872), .A2(G1991), .ZN(n980) );
  OR2_X1 U791 ( .A1(n974), .A2(n980), .ZN(n716) );
  NAND2_X1 U792 ( .A1(n716), .A2(n753), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n751), .A2(n743), .ZN(n717) );
  XOR2_X1 U794 ( .A(KEYINPUT87), .B(n717), .Z(n735) );
  OR2_X1 U795 ( .A1(n718), .A2(n735), .ZN(n719) );
  NOR2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n737) );
  INV_X1 U797 ( .A(n721), .ZN(n729) );
  NOR2_X1 U798 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U799 ( .A1(G8), .A2(n722), .ZN(n727) );
  NOR2_X1 U800 ( .A1(G1981), .A2(G305), .ZN(n723) );
  XOR2_X1 U801 ( .A(n723), .B(KEYINPUT88), .Z(n724) );
  XNOR2_X1 U802 ( .A(KEYINPUT24), .B(n724), .ZN(n725) );
  NOR2_X1 U803 ( .A1(n730), .A2(n725), .ZN(n731) );
  INV_X1 U804 ( .A(n731), .ZN(n726) );
  AND2_X1 U805 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n733) );
  OR2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n736) );
  OR2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U811 ( .A(n738), .B(KEYINPUT96), .ZN(n740) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n932) );
  NAND2_X1 U813 ( .A1(n932), .A2(n753), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n756) );
  NAND2_X1 U815 ( .A1(n741), .A2(n873), .ZN(n985) );
  XOR2_X1 U816 ( .A(KEYINPUT39), .B(KEYINPUT98), .Z(n749) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n844), .ZN(n742) );
  XOR2_X1 U818 ( .A(KEYINPUT97), .B(n742), .Z(n971) );
  INV_X1 U819 ( .A(n743), .ZN(n746) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n872), .ZN(n976) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n744) );
  NOR2_X1 U822 ( .A1(n976), .A2(n744), .ZN(n745) );
  NOR2_X1 U823 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U824 ( .A1(n971), .A2(n747), .ZN(n748) );
  XOR2_X1 U825 ( .A(n749), .B(n748), .Z(n750) );
  NAND2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n985), .A2(n752), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U831 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n825) );
  NAND2_X1 U837 ( .A1(n825), .A2(G567), .ZN(n760) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n760), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n766) );
  OR2_X1 U840 ( .A1(n936), .A2(n766), .ZN(n761) );
  XNOR2_X1 U841 ( .A(KEYINPUT72), .B(n761), .ZN(G153) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n763) );
  INV_X1 U843 ( .A(G868), .ZN(n806) );
  NAND2_X1 U844 ( .A1(n921), .A2(n806), .ZN(n762) );
  NAND2_X1 U845 ( .A1(n763), .A2(n762), .ZN(G284) );
  INV_X1 U846 ( .A(n924), .ZN(G299) );
  NOR2_X1 U847 ( .A1(G286), .A2(n806), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n766), .A2(G559), .ZN(n767) );
  INV_X1 U851 ( .A(n921), .ZN(n783) );
  NAND2_X1 U852 ( .A1(n767), .A2(n783), .ZN(n768) );
  XNOR2_X1 U853 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U854 ( .A1(G868), .A2(n936), .ZN(n771) );
  NAND2_X1 U855 ( .A1(G868), .A2(n783), .ZN(n769) );
  NOR2_X1 U856 ( .A1(G559), .A2(n769), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G123), .A2(n857), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT18), .ZN(n773) );
  XNOR2_X1 U860 ( .A(KEYINPUT74), .B(n773), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G111), .A2(n858), .ZN(n774) );
  XOR2_X1 U862 ( .A(KEYINPUT75), .B(n774), .Z(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U864 ( .A1(G99), .A2(n862), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G135), .A2(n865), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n973) );
  XNOR2_X1 U868 ( .A(n973), .B(G2096), .ZN(n782) );
  INV_X1 U869 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U871 ( .A1(n783), .A2(G559), .ZN(n803) );
  XNOR2_X1 U872 ( .A(n936), .B(n803), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n784), .A2(G860), .ZN(n795) );
  NAND2_X1 U874 ( .A1(G67), .A2(n785), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G93), .A2(n786), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G80), .A2(n789), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G55), .A2(n790), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n807) );
  XOR2_X1 U881 ( .A(n795), .B(n807), .Z(G145) );
  XNOR2_X1 U882 ( .A(n924), .B(G288), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(n807), .ZN(n801) );
  XNOR2_X1 U884 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U885 ( .A(G290), .B(G166), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U887 ( .A(G305), .B(n799), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n801), .B(n800), .ZN(n802) );
  XOR2_X1 U889 ( .A(n802), .B(n936), .Z(n829) );
  XOR2_X1 U890 ( .A(n829), .B(n803), .Z(n804) );
  NAND2_X1 U891 ( .A1(G868), .A2(n804), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n805), .B(KEYINPUT80), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2084), .A2(G2078), .ZN(n810) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XOR2_X1 U900 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  XNOR2_X1 U901 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U902 ( .A1(G69), .A2(G120), .ZN(n814) );
  NOR2_X1 U903 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U904 ( .A1(G108), .A2(n815), .ZN(n919) );
  NAND2_X1 U905 ( .A1(G567), .A2(n919), .ZN(n816) );
  XNOR2_X1 U906 ( .A(n816), .B(KEYINPUT81), .ZN(n821) );
  NOR2_X1 U907 ( .A1(G219), .A2(G220), .ZN(n817) );
  XNOR2_X1 U908 ( .A(KEYINPUT22), .B(n817), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(G96), .ZN(n819) );
  OR2_X1 U910 ( .A1(G218), .A2(n819), .ZN(n920) );
  AND2_X1 U911 ( .A1(G2106), .A2(n920), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n821), .A2(n820), .ZN(G319) );
  NAND2_X1 U913 ( .A1(G661), .A2(G483), .ZN(n823) );
  INV_X1 U914 ( .A(G319), .ZN(n822) );
  NOR2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(KEYINPUT82), .ZN(n828) );
  NAND2_X1 U917 ( .A1(G36), .A2(n828), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U923 ( .A(G96), .B(KEYINPUT100), .Z(G221) );
  XNOR2_X1 U924 ( .A(G286), .B(n921), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(G301), .ZN(n832) );
  NOR2_X1 U927 ( .A1(G37), .A2(n832), .ZN(G397) );
  NAND2_X1 U928 ( .A1(G124), .A2(n857), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT108), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n834), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U931 ( .A1(G100), .A2(n862), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n840) );
  NAND2_X1 U933 ( .A1(G112), .A2(n858), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G136), .A2(n865), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G162) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n843), .B(n973), .Z(n846) );
  XOR2_X1 U941 ( .A(n844), .B(G162), .Z(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n871) );
  NAND2_X1 U943 ( .A1(G106), .A2(n862), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G142), .A2(n865), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT45), .ZN(n856) );
  NAND2_X1 U947 ( .A1(n858), .A2(G118), .ZN(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT110), .B(n850), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n857), .A2(G130), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT109), .B(n851), .Z(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT111), .B(n854), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n869) );
  NAND2_X1 U954 ( .A1(G127), .A2(n857), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G115), .A2(n858), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n861), .B(KEYINPUT47), .ZN(n864) );
  NAND2_X1 U958 ( .A1(G103), .A2(n862), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U960 ( .A1(G139), .A2(n865), .ZN(n866) );
  XNOR2_X1 U961 ( .A(KEYINPUT113), .B(n866), .ZN(n867) );
  NOR2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n988) );
  XNOR2_X1 U963 ( .A(n869), .B(n988), .ZN(n870) );
  XNOR2_X1 U964 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U965 ( .A(n873), .B(n872), .Z(n874) );
  XNOR2_X1 U966 ( .A(n875), .B(n874), .ZN(n877) );
  XOR2_X1 U967 ( .A(G160), .B(G164), .Z(n876) );
  XNOR2_X1 U968 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U969 ( .A1(G37), .A2(n878), .ZN(G395) );
  XNOR2_X1 U970 ( .A(G1348), .B(G2454), .ZN(n879) );
  XNOR2_X1 U971 ( .A(n879), .B(G2430), .ZN(n880) );
  XNOR2_X1 U972 ( .A(n880), .B(G1341), .ZN(n886) );
  XOR2_X1 U973 ( .A(G2443), .B(G2427), .Z(n882) );
  XNOR2_X1 U974 ( .A(G2438), .B(G2446), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U976 ( .A(G2451), .B(G2435), .Z(n883) );
  XNOR2_X1 U977 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U978 ( .A(n886), .B(n885), .ZN(n887) );
  NAND2_X1 U979 ( .A1(n887), .A2(G14), .ZN(n888) );
  XNOR2_X1 U980 ( .A(KEYINPUT99), .B(n888), .ZN(G401) );
  XOR2_X1 U981 ( .A(G1961), .B(G1986), .Z(n890) );
  XNOR2_X1 U982 ( .A(G1996), .B(G1991), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n890), .B(n889), .ZN(n902) );
  XOR2_X1 U984 ( .A(G1976), .B(G1981), .Z(n892) );
  XNOR2_X1 U985 ( .A(G1956), .B(G1971), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U987 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n894) );
  XNOR2_X1 U988 ( .A(G1966), .B(KEYINPUT41), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U991 ( .A(G2474), .B(KEYINPUT107), .Z(n898) );
  XNOR2_X1 U992 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(G229) );
  XOR2_X1 U996 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n904) );
  XNOR2_X1 U997 ( .A(KEYINPUT101), .B(G2678), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U999 ( .A(KEYINPUT42), .B(G2090), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G2067), .B(G2072), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G2096), .B(G2100), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1005 ( .A(G2084), .B(G2078), .Z(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(G227) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n913) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n914), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n915), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G397), .A2(G395), .ZN(n916) );
  XOR2_X1 U1012 ( .A(KEYINPUT115), .B(n916), .Z(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  XOR2_X1 U1014 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1016 ( .A(G120), .ZN(G236) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1019 ( .A(G325), .ZN(G261) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(KEYINPUT56), .B(G16), .ZN(n947) );
  XNOR2_X1 U1022 ( .A(G301), .B(G1961), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n921), .B(G1348), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(G166), .B(G1971), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n924), .B(G1956), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1031 ( .A(KEYINPUT123), .B(n933), .Z(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(G1341), .B(n936), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT57), .ZN(n943) );
  XOR2_X1 U1038 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n942) );
  XNOR2_X1 U1039 ( .A(n943), .B(n942), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(KEYINPUT124), .B(n948), .ZN(n1001) );
  XOR2_X1 U1043 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n966) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n961) );
  XOR2_X1 U1045 ( .A(G25), .B(G1991), .Z(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G27), .B(n952), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n966), .B(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G29), .B(KEYINPUT120), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n999) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1066 ( .A(KEYINPUT51), .B(n972), .Z(n982) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n978) );
  XOR2_X1 U1068 ( .A(G160), .B(G2084), .Z(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1075 ( .A(KEYINPUT117), .B(n987), .Z(n993) );
  XOR2_X1 U1076 ( .A(G2072), .B(n988), .Z(n990) );
  XOR2_X1 U1077 ( .A(G164), .B(G2078), .Z(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT50), .B(n991), .Z(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1081 ( .A(KEYINPUT52), .B(n994), .Z(n995) );
  NOR2_X1 U1082 ( .A1(KEYINPUT55), .A2(n995), .ZN(n997) );
  INV_X1 U1083 ( .A(G29), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1029) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(n1002), .B(G4), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(G1348), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1010), .B(KEYINPUT60), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G1986), .B(KEYINPUT127), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1016), .B(G24), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1019), .Z(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G5), .B(G1961), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1024), .ZN(n1026) );
  INV_X1 U1111 ( .A(G16), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(n1030), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

