

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n683), .A2(n577), .ZN(n693) );
  AND2_X1 U551 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U552 ( .A(n757), .ZN(n730) );
  XNOR2_X1 U553 ( .A(KEYINPUT68), .B(n579), .ZN(n690) );
  XNOR2_X1 U554 ( .A(n576), .B(KEYINPUT86), .ZN(G164) );
  XNOR2_X2 U555 ( .A(n565), .B(n563), .ZN(n610) );
  NOR2_X2 U556 ( .A1(n764), .A2(n763), .ZN(n765) );
  BUF_X2 U557 ( .A(n587), .Z(n517) );
  OR2_X1 U558 ( .A1(n782), .A2(n781), .ZN(n786) );
  NOR2_X1 U559 ( .A1(n772), .A2(G1966), .ZN(n768) );
  XNOR2_X1 U560 ( .A(n758), .B(KEYINPUT91), .ZN(n797) );
  AND2_X1 U561 ( .A1(G160), .A2(G40), .ZN(n727) );
  BUF_X1 U562 ( .A(n610), .Z(n588) );
  NOR2_X2 U563 ( .A1(G2105), .A2(n573), .ZN(n587) );
  XNOR2_X1 U564 ( .A(KEYINPUT66), .B(KEYINPUT17), .ZN(n565) );
  XNOR2_X1 U565 ( .A(n765), .B(KEYINPUT31), .ZN(n771) );
  INV_X1 U566 ( .A(KEYINPUT40), .ZN(n537) );
  NOR2_X1 U567 ( .A1(n527), .A2(G299), .ZN(n747) );
  XNOR2_X1 U568 ( .A(KEYINPUT32), .B(KEYINPUT99), .ZN(n787) );
  NAND2_X1 U569 ( .A1(n543), .A2(n524), .ZN(n542) );
  NAND2_X1 U570 ( .A1(n525), .A2(n549), .ZN(n543) );
  NAND2_X1 U571 ( .A1(n796), .A2(n518), .ZN(n540) );
  NOR2_X1 U572 ( .A1(n538), .A2(n537), .ZN(n536) );
  NAND2_X1 U573 ( .A1(n534), .A2(n533), .ZN(n532) );
  NAND2_X1 U574 ( .A1(n863), .A2(n526), .ZN(n533) );
  NAND2_X1 U575 ( .A1(n535), .A2(n537), .ZN(n534) );
  INV_X1 U576 ( .A(KEYINPUT23), .ZN(n615) );
  NAND2_X1 U577 ( .A1(n745), .A2(n744), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n558), .B(n557), .ZN(n782) );
  INV_X1 U579 ( .A(KEYINPUT96), .ZN(n557) );
  NOR2_X1 U580 ( .A1(n546), .A2(KEYINPUT103), .ZN(n545) );
  INV_X1 U581 ( .A(n522), .ZN(n546) );
  NOR2_X1 U582 ( .A1(n768), .A2(n523), .ZN(n769) );
  NAND2_X1 U583 ( .A1(n757), .A2(G8), .ZN(n758) );
  NOR2_X1 U584 ( .A1(G164), .A2(G1384), .ZN(n817) );
  INV_X1 U585 ( .A(n863), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n627), .B(KEYINPUT71), .ZN(n628) );
  NAND2_X1 U587 ( .A1(n573), .A2(n564), .ZN(n563) );
  INV_X1 U588 ( .A(G2105), .ZN(n564) );
  NOR2_X1 U589 ( .A1(G651), .A2(n683), .ZN(n697) );
  NAND2_X1 U590 ( .A1(n530), .A2(n519), .ZN(n529) );
  INV_X1 U591 ( .A(KEYINPUT64), .ZN(n560) );
  AND2_X1 U592 ( .A1(n549), .A2(KEYINPUT103), .ZN(n518) );
  INV_X1 U593 ( .A(n797), .ZN(n772) );
  INV_X1 U594 ( .A(n797), .ZN(n549) );
  AND2_X1 U595 ( .A1(n863), .A2(n537), .ZN(n519) );
  XNOR2_X1 U596 ( .A(KEYINPUT93), .B(n756), .ZN(n520) );
  AND2_X1 U597 ( .A1(n555), .A2(n554), .ZN(n521) );
  OR2_X1 U598 ( .A1(G2090), .A2(n791), .ZN(n522) );
  AND2_X1 U599 ( .A1(n767), .A2(G8), .ZN(n523) );
  OR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n524) );
  OR2_X1 U601 ( .A1(n522), .A2(n548), .ZN(n525) );
  INV_X1 U602 ( .A(KEYINPUT103), .ZN(n548) );
  OR2_X1 U603 ( .A1(n851), .A2(KEYINPUT40), .ZN(n526) );
  NAND2_X1 U604 ( .A1(n527), .A2(G299), .ZN(n750) );
  AND2_X1 U605 ( .A1(n528), .A2(n532), .ZN(n531) );
  NAND2_X1 U606 ( .A1(n539), .A2(n536), .ZN(n528) );
  XNOR2_X1 U607 ( .A(n850), .B(n849), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n531), .A2(n529), .ZN(G329) );
  INV_X1 U609 ( .A(n539), .ZN(n530) );
  INV_X1 U610 ( .A(n851), .ZN(n538) );
  NAND2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n547) );
  AND2_X1 U612 ( .A1(n544), .A2(n542), .ZN(n541) );
  NAND2_X1 U613 ( .A1(n550), .A2(n545), .ZN(n544) );
  NAND2_X1 U614 ( .A1(n809), .A2(n547), .ZN(n810) );
  INV_X1 U615 ( .A(n796), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n521), .A2(n551), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n551) );
  INV_X1 U618 ( .A(n753), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n752), .A2(n556), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n752), .A2(n556), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n753), .A2(n556), .ZN(n555) );
  INV_X1 U622 ( .A(KEYINPUT29), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n559), .A2(n520), .ZN(n558) );
  XNOR2_X2 U624 ( .A(n561), .B(n560), .ZN(G160) );
  NAND2_X1 U625 ( .A1(n562), .A2(n619), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n614), .B(KEYINPUT67), .ZN(n562) );
  NOR2_X2 U627 ( .A1(n790), .A2(n789), .ZN(n796) );
  AND2_X1 U628 ( .A1(n770), .A2(n769), .ZN(n790) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n622), .Z(n566) );
  INV_X1 U630 ( .A(KEYINPUT26), .ZN(n731) );
  INV_X1 U631 ( .A(KEYINPUT27), .ZN(n742) );
  INV_X1 U632 ( .A(KEYINPUT95), .ZN(n746) );
  INV_X1 U633 ( .A(KEYINPUT13), .ZN(n627) );
  INV_X1 U634 ( .A(KEYINPUT105), .ZN(n849) );
  INV_X1 U635 ( .A(G651), .ZN(n577) );
  XNOR2_X1 U636 ( .A(n629), .B(n628), .ZN(n630) );
  AND2_X1 U637 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U638 ( .A1(G2105), .A2(G2104), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT65), .ZN(n611) );
  NAND2_X1 U640 ( .A1(G114), .A2(n611), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G138), .A2(n610), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n572) );
  INV_X1 U643 ( .A(G2104), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G102), .A2(n587), .ZN(n570) );
  XNOR2_X1 U645 ( .A(KEYINPUT85), .B(n570), .ZN(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n575) );
  AND2_X1 U647 ( .A1(n573), .A2(G2105), .ZN(n916) );
  NAND2_X1 U648 ( .A1(n916), .A2(G126), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT0), .B(G543), .Z(n683) );
  NAND2_X1 U650 ( .A1(n693), .A2(G78), .ZN(n581) );
  NOR2_X1 U651 ( .A1(G543), .A2(n577), .ZN(n578) );
  XOR2_X1 U652 ( .A(KEYINPUT1), .B(n578), .Z(n579) );
  NAND2_X1 U653 ( .A1(G65), .A2(n690), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n585) );
  NOR2_X1 U655 ( .A1(G651), .A2(G543), .ZN(n689) );
  NAND2_X1 U656 ( .A1(G91), .A2(n689), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G53), .A2(n697), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U659 ( .A1(n585), .A2(n584), .ZN(G299) );
  AND2_X1 U660 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U661 ( .A(n611), .Z(n915) );
  NAND2_X1 U662 ( .A1(G111), .A2(n915), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT76), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G99), .A2(n517), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G135), .A2(n588), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n916), .A2(G123), .ZN(n591) );
  XOR2_X1 U668 ( .A(KEYINPUT18), .B(n591), .Z(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n1030) );
  XNOR2_X1 U671 ( .A(G2096), .B(n1030), .ZN(n596) );
  OR2_X1 U672 ( .A1(G2100), .A2(n596), .ZN(G156) );
  INV_X1 U673 ( .A(G57), .ZN(G237) );
  INV_X1 U674 ( .A(G132), .ZN(G219) );
  INV_X1 U675 ( .A(G82), .ZN(G220) );
  NAND2_X1 U676 ( .A1(n693), .A2(G76), .ZN(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT73), .B(n597), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n689), .A2(G89), .ZN(n598) );
  XOR2_X1 U679 ( .A(n598), .B(KEYINPUT4), .Z(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U681 ( .A(KEYINPUT5), .B(n601), .Z(n602) );
  XNOR2_X1 U682 ( .A(KEYINPUT74), .B(n602), .ZN(n608) );
  XNOR2_X1 U683 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n697), .A2(G51), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G63), .A2(n690), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U690 ( .A1(n610), .A2(G137), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G113), .A2(n611), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G125), .A2(n916), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G101), .A2(n517), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(n615), .ZN(n617) );
  XOR2_X1 U696 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U697 ( .A1(G7), .A2(G661), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U699 ( .A(G223), .ZN(n864) );
  NAND2_X1 U700 ( .A1(n864), .A2(G567), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT11), .B(n621), .Z(G234) );
  NAND2_X1 U702 ( .A1(G56), .A2(n690), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n689), .A2(G81), .ZN(n623) );
  XOR2_X1 U704 ( .A(KEYINPUT12), .B(n623), .Z(n626) );
  NAND2_X1 U705 ( .A1(n693), .A2(G68), .ZN(n624) );
  XOR2_X1 U706 ( .A(n624), .B(KEYINPUT70), .Z(n625) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n566), .A2(n630), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n697), .A2(G43), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n1008) );
  INV_X1 U711 ( .A(G860), .ZN(n653) );
  OR2_X1 U712 ( .A1(n1008), .A2(n653), .ZN(G153) );
  NAND2_X1 U713 ( .A1(n690), .A2(G64), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n633), .B(KEYINPUT69), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G77), .A2(n693), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G90), .A2(n689), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U718 ( .A(KEYINPUT9), .B(n636), .Z(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n697), .A2(G52), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(G301) );
  NAND2_X1 U722 ( .A1(G868), .A2(G301), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n689), .A2(G92), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G66), .A2(n690), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G79), .A2(n693), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G54), .A2(n697), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U729 ( .A(KEYINPUT72), .B(n645), .ZN(n646) );
  NOR2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT15), .ZN(n739) );
  INV_X1 U732 ( .A(G868), .ZN(n708) );
  NAND2_X1 U733 ( .A1(n739), .A2(n708), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G284) );
  NOR2_X1 U735 ( .A1(G286), .A2(n708), .ZN(n652) );
  NOR2_X1 U736 ( .A1(G868), .A2(G299), .ZN(n651) );
  NOR2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G297) );
  NAND2_X1 U738 ( .A1(n653), .A2(G559), .ZN(n654) );
  INV_X1 U739 ( .A(n739), .ZN(n1001) );
  NAND2_X1 U740 ( .A1(n654), .A2(n1001), .ZN(n655) );
  XNOR2_X1 U741 ( .A(n655), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U742 ( .A1(G868), .A2(n1008), .ZN(n658) );
  NAND2_X1 U743 ( .A1(G868), .A2(n1001), .ZN(n656) );
  NOR2_X1 U744 ( .A1(G559), .A2(n656), .ZN(n657) );
  NOR2_X1 U745 ( .A1(n658), .A2(n657), .ZN(G282) );
  NAND2_X1 U746 ( .A1(G559), .A2(n1001), .ZN(n659) );
  XNOR2_X1 U747 ( .A(n659), .B(n1008), .ZN(n706) );
  NOR2_X1 U748 ( .A1(n706), .A2(G860), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n689), .A2(G93), .ZN(n660) );
  XOR2_X1 U750 ( .A(KEYINPUT77), .B(n660), .Z(n662) );
  NAND2_X1 U751 ( .A1(n693), .A2(G80), .ZN(n661) );
  NAND2_X1 U752 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U753 ( .A(KEYINPUT78), .B(n663), .Z(n665) );
  NAND2_X1 U754 ( .A1(G67), .A2(n690), .ZN(n664) );
  NAND2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U756 ( .A1(G55), .A2(n697), .ZN(n666) );
  XNOR2_X1 U757 ( .A(KEYINPUT79), .B(n666), .ZN(n667) );
  OR2_X1 U758 ( .A1(n668), .A2(n667), .ZN(n709) );
  XOR2_X1 U759 ( .A(n669), .B(n709), .Z(G145) );
  AND2_X1 U760 ( .A1(G60), .A2(n690), .ZN(n673) );
  NAND2_X1 U761 ( .A1(G72), .A2(n693), .ZN(n671) );
  NAND2_X1 U762 ( .A1(G85), .A2(n689), .ZN(n670) );
  NAND2_X1 U763 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U764 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U765 ( .A1(n697), .A2(G47), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n675), .A2(n674), .ZN(G290) );
  NAND2_X1 U767 ( .A1(G75), .A2(n693), .ZN(n677) );
  NAND2_X1 U768 ( .A1(G88), .A2(n689), .ZN(n676) );
  NAND2_X1 U769 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n697), .A2(G50), .ZN(n678) );
  XOR2_X1 U771 ( .A(KEYINPUT80), .B(n678), .Z(n679) );
  NOR2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U773 ( .A1(G62), .A2(n690), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n682), .A2(n681), .ZN(G303) );
  INV_X1 U775 ( .A(G303), .ZN(G166) );
  NAND2_X1 U776 ( .A1(G87), .A2(n683), .ZN(n685) );
  NAND2_X1 U777 ( .A1(G74), .A2(G651), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n690), .A2(n686), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n697), .A2(G49), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(G288) );
  NAND2_X1 U782 ( .A1(n689), .A2(G86), .ZN(n692) );
  NAND2_X1 U783 ( .A1(G61), .A2(n690), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n693), .A2(G73), .ZN(n694) );
  XOR2_X1 U786 ( .A(KEYINPUT2), .B(n694), .Z(n695) );
  NOR2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n697), .A2(G48), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(G305) );
  XNOR2_X1 U790 ( .A(G290), .B(G299), .ZN(n705) );
  XNOR2_X1 U791 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n701) );
  XOR2_X1 U792 ( .A(G288), .B(n709), .Z(n700) );
  XNOR2_X1 U793 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U794 ( .A(G166), .B(n702), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(G305), .ZN(n704) );
  XNOR2_X1 U796 ( .A(n705), .B(n704), .ZN(n934) );
  XNOR2_X1 U797 ( .A(n706), .B(n934), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n707), .A2(G868), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(G295) );
  NAND2_X1 U801 ( .A1(G2084), .A2(G2078), .ZN(n712) );
  XOR2_X1 U802 ( .A(KEYINPUT20), .B(n712), .Z(n713) );
  NAND2_X1 U803 ( .A1(G2090), .A2(n713), .ZN(n714) );
  XNOR2_X1 U804 ( .A(KEYINPUT21), .B(n714), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n715), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT82), .B(n716), .ZN(G158) );
  XOR2_X1 U807 ( .A(KEYINPUT83), .B(G44), .Z(n717) );
  XNOR2_X1 U808 ( .A(KEYINPUT3), .B(n717), .ZN(G218) );
  NOR2_X1 U809 ( .A1(G220), .A2(G219), .ZN(n718) );
  XOR2_X1 U810 ( .A(KEYINPUT22), .B(n718), .Z(n719) );
  NOR2_X1 U811 ( .A1(G218), .A2(n719), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT84), .B(n720), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n721), .A2(G96), .ZN(n871) );
  NAND2_X1 U814 ( .A1(n871), .A2(G2106), .ZN(n725) );
  NAND2_X1 U815 ( .A1(G120), .A2(G69), .ZN(n722) );
  NOR2_X1 U816 ( .A1(G237), .A2(n722), .ZN(n723) );
  NAND2_X1 U817 ( .A1(G108), .A2(n723), .ZN(n872) );
  NAND2_X1 U818 ( .A1(n872), .A2(G567), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n873) );
  NAND2_X1 U820 ( .A1(G661), .A2(G483), .ZN(n726) );
  NOR2_X1 U821 ( .A1(n873), .A2(n726), .ZN(n868) );
  NAND2_X1 U822 ( .A1(n868), .A2(G36), .ZN(G176) );
  INV_X1 U823 ( .A(G301), .ZN(G171) );
  NAND2_X2 U824 ( .A1(n727), .A2(n817), .ZN(n757) );
  NAND2_X1 U825 ( .A1(n730), .A2(G2067), .ZN(n729) );
  NAND2_X1 U826 ( .A1(G1348), .A2(n757), .ZN(n728) );
  NAND2_X1 U827 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n738), .A2(n739), .ZN(n737) );
  AND2_X1 U829 ( .A1(n730), .A2(G1996), .ZN(n732) );
  XNOR2_X1 U830 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U831 ( .A1(n757), .A2(G1341), .ZN(n733) );
  NAND2_X1 U832 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U833 ( .A1(n735), .A2(n1008), .ZN(n736) );
  NOR2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X2 U836 ( .A1(n741), .A2(n740), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n730), .A2(G2072), .ZN(n743) );
  XNOR2_X1 U838 ( .A(n743), .B(n742), .ZN(n745) );
  NAND2_X1 U839 ( .A1(G1956), .A2(n757), .ZN(n744) );
  XNOR2_X1 U840 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X2 U841 ( .A1(n749), .A2(n748), .ZN(n753) );
  XOR2_X1 U842 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U844 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NOR2_X1 U845 ( .A1(n757), .A2(n958), .ZN(n755) );
  AND2_X1 U846 ( .A1(n757), .A2(G1961), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n762) );
  AND2_X1 U848 ( .A1(G171), .A2(n762), .ZN(n756) );
  NOR2_X1 U849 ( .A1(G2084), .A2(n757), .ZN(n767) );
  NOR2_X1 U850 ( .A1(n768), .A2(n767), .ZN(n759) );
  NAND2_X1 U851 ( .A1(G8), .A2(n759), .ZN(n760) );
  XNOR2_X1 U852 ( .A(KEYINPUT30), .B(n760), .ZN(n761) );
  NOR2_X1 U853 ( .A1(G168), .A2(n761), .ZN(n764) );
  NOR2_X1 U854 ( .A1(G171), .A2(n762), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n782), .A2(n771), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT97), .ZN(n770) );
  INV_X1 U857 ( .A(n771), .ZN(n780) );
  INV_X1 U858 ( .A(G8), .ZN(n778) );
  NOR2_X1 U859 ( .A1(G1971), .A2(n549), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n757), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n775), .A2(G303), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n776), .B(KEYINPUT98), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n784) );
  INV_X1 U865 ( .A(n784), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U867 ( .A1(G286), .A2(G8), .ZN(n783) );
  OR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n786), .A2(n785), .ZN(n788) );
  XNOR2_X1 U870 ( .A(n788), .B(n787), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G166), .A2(G8), .ZN(n791) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  NOR2_X1 U873 ( .A1(G1971), .A2(G303), .ZN(n792) );
  XNOR2_X1 U874 ( .A(KEYINPUT100), .B(n792), .ZN(n793) );
  NOR2_X1 U875 ( .A1(n1012), .A2(n793), .ZN(n794) );
  XNOR2_X1 U876 ( .A(n794), .B(KEYINPUT101), .ZN(n795) );
  NOR2_X1 U877 ( .A1(n796), .A2(n795), .ZN(n805) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NAND2_X1 U879 ( .A1(n1013), .A2(n797), .ZN(n803) );
  NAND2_X1 U880 ( .A1(n1012), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U881 ( .A1(n798), .A2(n549), .ZN(n801) );
  XOR2_X1 U882 ( .A(G1981), .B(KEYINPUT102), .Z(n799) );
  XNOR2_X1 U883 ( .A(G305), .B(n799), .ZN(n1003) );
  INV_X1 U884 ( .A(n1003), .ZN(n800) );
  NOR2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n806) );
  INV_X1 U886 ( .A(n806), .ZN(n802) );
  OR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U888 ( .A1(n805), .A2(n804), .ZN(n808) );
  AND2_X1 U889 ( .A1(n806), .A2(KEYINPUT33), .ZN(n807) );
  NOR2_X1 U890 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U891 ( .A(n810), .B(KEYINPUT104), .ZN(n815) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U893 ( .A(n811), .B(KEYINPUT24), .Z(n812) );
  XNOR2_X1 U894 ( .A(KEYINPUT92), .B(n812), .ZN(n813) );
  NOR2_X1 U895 ( .A1(n549), .A2(n813), .ZN(n814) );
  NOR2_X1 U896 ( .A1(n815), .A2(n814), .ZN(n848) );
  NAND2_X1 U897 ( .A1(G40), .A2(G160), .ZN(n816) );
  NOR2_X1 U898 ( .A1(n817), .A2(n816), .ZN(n861) );
  NAND2_X1 U899 ( .A1(n517), .A2(G104), .ZN(n818) );
  XOR2_X1 U900 ( .A(KEYINPUT87), .B(n818), .Z(n820) );
  NAND2_X1 U901 ( .A1(G140), .A2(n588), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U903 ( .A(KEYINPUT34), .B(n821), .ZN(n826) );
  NAND2_X1 U904 ( .A1(G116), .A2(n915), .ZN(n823) );
  NAND2_X1 U905 ( .A1(G128), .A2(n916), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U907 ( .A(KEYINPUT35), .B(n824), .Z(n825) );
  NOR2_X1 U908 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n827), .ZN(n901) );
  XNOR2_X1 U910 ( .A(G2067), .B(KEYINPUT37), .ZN(n858) );
  NOR2_X1 U911 ( .A1(n901), .A2(n858), .ZN(n1040) );
  NAND2_X1 U912 ( .A1(n861), .A2(n1040), .ZN(n856) );
  NAND2_X1 U913 ( .A1(n916), .A2(G119), .ZN(n834) );
  NAND2_X1 U914 ( .A1(G107), .A2(n915), .ZN(n829) );
  NAND2_X1 U915 ( .A1(G131), .A2(n588), .ZN(n828) );
  NAND2_X1 U916 ( .A1(n829), .A2(n828), .ZN(n832) );
  NAND2_X1 U917 ( .A1(n517), .A2(G95), .ZN(n830) );
  XOR2_X1 U918 ( .A(KEYINPUT88), .B(n830), .Z(n831) );
  NOR2_X1 U919 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U921 ( .A(KEYINPUT89), .B(n835), .Z(n903) );
  NAND2_X1 U922 ( .A1(G1991), .A2(n903), .ZN(n836) );
  XNOR2_X1 U923 ( .A(n836), .B(KEYINPUT90), .ZN(n845) );
  NAND2_X1 U924 ( .A1(G117), .A2(n915), .ZN(n838) );
  NAND2_X1 U925 ( .A1(G141), .A2(n588), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n838), .A2(n837), .ZN(n841) );
  NAND2_X1 U927 ( .A1(n517), .A2(G105), .ZN(n839) );
  XOR2_X1 U928 ( .A(KEYINPUT38), .B(n839), .Z(n840) );
  NOR2_X1 U929 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U930 ( .A1(n916), .A2(G129), .ZN(n842) );
  NAND2_X1 U931 ( .A1(n843), .A2(n842), .ZN(n927) );
  NAND2_X1 U932 ( .A1(G1996), .A2(n927), .ZN(n844) );
  NAND2_X1 U933 ( .A1(n845), .A2(n844), .ZN(n1029) );
  NAND2_X1 U934 ( .A1(n861), .A2(n1029), .ZN(n846) );
  NAND2_X1 U935 ( .A1(n856), .A2(n846), .ZN(n847) );
  NOR2_X1 U936 ( .A1(n848), .A2(n847), .ZN(n850) );
  XNOR2_X1 U937 ( .A(G1986), .B(G290), .ZN(n1020) );
  NAND2_X1 U938 ( .A1(n1020), .A2(n861), .ZN(n851) );
  NOR2_X1 U939 ( .A1(G1996), .A2(n927), .ZN(n1037) );
  NOR2_X1 U940 ( .A1(G1986), .A2(G290), .ZN(n852) );
  NOR2_X1 U941 ( .A1(G1991), .A2(n903), .ZN(n1033) );
  NOR2_X1 U942 ( .A1(n852), .A2(n1033), .ZN(n853) );
  NOR2_X1 U943 ( .A1(n1029), .A2(n853), .ZN(n854) );
  NOR2_X1 U944 ( .A1(n1037), .A2(n854), .ZN(n855) );
  XNOR2_X1 U945 ( .A(n855), .B(KEYINPUT39), .ZN(n857) );
  NAND2_X1 U946 ( .A1(n857), .A2(n856), .ZN(n859) );
  NAND2_X1 U947 ( .A1(n901), .A2(n858), .ZN(n1031) );
  NAND2_X1 U948 ( .A1(n859), .A2(n1031), .ZN(n860) );
  NAND2_X1 U949 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U950 ( .A(KEYINPUT106), .B(n862), .ZN(n863) );
  NAND2_X1 U951 ( .A1(G2106), .A2(n864), .ZN(G217) );
  INV_X1 U952 ( .A(G661), .ZN(n866) );
  NAND2_X1 U953 ( .A1(G2), .A2(G15), .ZN(n865) );
  NOR2_X1 U954 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U955 ( .A(KEYINPUT108), .B(n867), .Z(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n869) );
  NAND2_X1 U957 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(n870), .Z(G188) );
  XOR2_X1 U959 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U961 ( .A(G120), .ZN(G236) );
  INV_X1 U962 ( .A(G96), .ZN(G221) );
  NOR2_X1 U963 ( .A1(n872), .A2(n871), .ZN(G325) );
  INV_X1 U964 ( .A(G325), .ZN(G261) );
  INV_X1 U965 ( .A(n873), .ZN(G319) );
  XOR2_X1 U966 ( .A(KEYINPUT42), .B(G2090), .Z(n875) );
  XNOR2_X1 U967 ( .A(G2084), .B(G2067), .ZN(n874) );
  XNOR2_X1 U968 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U969 ( .A(n876), .B(G2100), .Z(n878) );
  XNOR2_X1 U970 ( .A(G2078), .B(G2072), .ZN(n877) );
  XNOR2_X1 U971 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U972 ( .A(G2096), .B(KEYINPUT43), .Z(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(G2678), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U975 ( .A(n882), .B(n881), .Z(G227) );
  XOR2_X1 U976 ( .A(KEYINPUT41), .B(G1956), .Z(n884) );
  XNOR2_X1 U977 ( .A(G1976), .B(G1961), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U979 ( .A(n885), .B(KEYINPUT113), .Z(n887) );
  XNOR2_X1 U980 ( .A(G1996), .B(G1991), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U982 ( .A(G1971), .B(G1966), .Z(n889) );
  XNOR2_X1 U983 ( .A(G1986), .B(G1981), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(n891), .B(n890), .Z(n893) );
  XNOR2_X1 U986 ( .A(KEYINPUT112), .B(G2474), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(G229) );
  NAND2_X1 U988 ( .A1(G124), .A2(n916), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(KEYINPUT44), .ZN(n896) );
  NAND2_X1 U990 ( .A1(n915), .A2(G112), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G100), .A2(n517), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G136), .A2(n588), .ZN(n897) );
  NAND2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(G162) );
  XOR2_X1 U996 ( .A(G164), .B(n901), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n1030), .B(n904), .ZN(n914) );
  NAND2_X1 U999 ( .A1(G103), .A2(n517), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G139), .A2(n588), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n915), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n916), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(KEYINPUT47), .B(n909), .Z(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1007 ( .A(KEYINPUT116), .B(n912), .Z(n1041) );
  XNOR2_X1 U1008 ( .A(n1041), .B(G162), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n932) );
  NAND2_X1 U1010 ( .A1(G118), .A2(n915), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(G130), .A2(n916), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(KEYINPUT114), .B(n919), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(G106), .A2(n517), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(G142), .A2(n588), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1017 ( .A(n922), .B(KEYINPUT45), .Z(n923) );
  NOR2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1019 ( .A(KEYINPUT48), .B(n925), .Z(n926) );
  XNOR2_X1 U1020 ( .A(KEYINPUT46), .B(n926), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(n927), .B(KEYINPUT115), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(n929), .B(n928), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G160), .B(n930), .Z(n931) );
  XNOR2_X1 U1024 ( .A(n932), .B(n931), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n933), .ZN(G395) );
  XNOR2_X1 U1026 ( .A(n1008), .B(G286), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(n935), .B(n934), .ZN(n937) );
  XOR2_X1 U1028 ( .A(n1001), .B(G171), .Z(n936) );
  XNOR2_X1 U1029 ( .A(n937), .B(n936), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(G37), .A2(n938), .ZN(G397) );
  XOR2_X1 U1031 ( .A(G2430), .B(G2451), .Z(n940) );
  XNOR2_X1 U1032 ( .A(G2446), .B(G2427), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n940), .B(n939), .ZN(n947) );
  XOR2_X1 U1034 ( .A(G2438), .B(G2435), .Z(n942) );
  XNOR2_X1 U1035 ( .A(G2443), .B(KEYINPUT107), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n942), .B(n941), .ZN(n943) );
  XOR2_X1 U1037 ( .A(n943), .B(G2454), .Z(n945) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G1348), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n945), .B(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n947), .B(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G14), .ZN(n954) );
  NAND2_X1 U1042 ( .A1(G319), .A2(n954), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(G227), .A2(G229), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT49), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(G395), .A2(G397), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(G225) );
  INV_X1 U1048 ( .A(G225), .ZN(G308) );
  INV_X1 U1049 ( .A(G108), .ZN(G238) );
  INV_X1 U1050 ( .A(n954), .ZN(G401) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2072), .B(G33), .Z(n957) );
  NAND2_X1 U1055 ( .A1(n957), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G27), .B(n958), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G25), .B(G1991), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT53), .B(n966), .Z(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT54), .B(G34), .Z(n967) );
  XNOR2_X1 U1064 ( .A(G2084), .B(n967), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G35), .B(G2090), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n972), .Z(n973) );
  NOR2_X1 U1069 ( .A1(G29), .A2(n973), .ZN(n1057) );
  XNOR2_X1 U1070 ( .A(KEYINPUT121), .B(G16), .ZN(n1000) );
  XNOR2_X1 U1071 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(G1341), .B(G19), .ZN(n975) );
  NOR2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1077 ( .A(KEYINPUT123), .B(G1956), .Z(n979) );
  XNOR2_X1 U1078 ( .A(G20), .B(n979), .ZN(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(KEYINPUT60), .B(n982), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G1961), .B(KEYINPUT122), .ZN(n983) );
  XNOR2_X1 U1082 ( .A(n983), .B(G5), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G1986), .B(G24), .ZN(n985) );
  XNOR2_X1 U1084 ( .A(G22), .B(G1971), .ZN(n984) );
  NOR2_X1 U1085 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1086 ( .A(G1976), .B(KEYINPUT125), .ZN(n986) );
  XNOR2_X1 U1087 ( .A(n986), .B(G23), .ZN(n987) );
  NAND2_X1 U1088 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n989), .ZN(n990) );
  NOR2_X1 U1090 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1092 ( .A(KEYINPUT124), .B(G1966), .ZN(n994) );
  XNOR2_X1 U1093 ( .A(G21), .B(n994), .ZN(n995) );
  NOR2_X1 U1094 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1095 ( .A(n997), .B(KEYINPUT126), .ZN(n998) );
  XNOR2_X1 U1096 ( .A(n998), .B(KEYINPUT61), .ZN(n999) );
  NAND2_X1 U1097 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  XNOR2_X1 U1098 ( .A(KEYINPUT56), .B(G16), .ZN(n1024) );
  XNOR2_X1 U1099 ( .A(G1348), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1100 ( .A(n1002), .B(KEYINPUT120), .ZN(n1007) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1102 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1103 ( .A(n1005), .B(KEYINPUT57), .ZN(n1006) );
  NAND2_X1 U1104 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1105 ( .A(G1341), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1106 ( .A1(n1010), .A2(n1009), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G166), .B(G1971), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G1956), .B(G299), .ZN(n1011) );
  NOR2_X1 U1109 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NAND2_X1 U1110 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1111 ( .A(G1961), .B(G301), .ZN(n1015) );
  NOR2_X1 U1112 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1113 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1114 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1115 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1116 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1117 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1118 ( .A(n1027), .B(KEYINPUT127), .ZN(n1055) );
  XOR2_X1 U1119 ( .A(G2084), .B(G160), .Z(n1028) );
  NOR2_X1 U1120 ( .A1(n1029), .A2(n1028), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1049) );
  XOR2_X1 U1124 ( .A(G2090), .B(G162), .Z(n1036) );
  NOR2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1126 ( .A(n1038), .B(KEYINPUT51), .ZN(n1039) );
  NOR2_X1 U1127 ( .A1(n1040), .A2(n1039), .ZN(n1047) );
  XOR2_X1 U1128 ( .A(G164), .B(G2078), .Z(n1043) );
  XNOR2_X1 U1129 ( .A(G2072), .B(n1041), .ZN(n1042) );
  NOR2_X1 U1130 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1131 ( .A(n1044), .B(KEYINPUT50), .Z(n1045) );
  XNOR2_X1 U1132 ( .A(KEYINPUT117), .B(n1045), .ZN(n1046) );
  NAND2_X1 U1133 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1134 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XOR2_X1 U1135 ( .A(KEYINPUT52), .B(n1050), .Z(n1051) );
  NOR2_X1 U1136 ( .A1(KEYINPUT55), .A2(n1051), .ZN(n1052) );
  XOR2_X1 U1137 ( .A(KEYINPUT118), .B(n1052), .Z(n1053) );
  NAND2_X1 U1138 ( .A1(n1053), .A2(G29), .ZN(n1054) );
  NAND2_X1 U1139 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NOR2_X1 U1140 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1141 ( .A1(n1058), .A2(G11), .ZN(n1059) );
  XOR2_X1 U1142 ( .A(KEYINPUT62), .B(n1059), .Z(G311) );
  INV_X1 U1143 ( .A(G311), .ZN(G150) );
endmodule

