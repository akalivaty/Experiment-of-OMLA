//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n187), .A2(new_n188), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT71), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT3), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n196), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n192), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n205), .B2(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n199), .A2(new_n197), .B1(new_n213), .B2(new_n196), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT72), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n200), .A2(new_n204), .A3(KEYINPUT72), .A4(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n210), .B(new_n211), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n200), .A2(new_n204), .A3(new_n215), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n217), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n210), .B1(new_n224), .B2(new_n211), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT76), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n211), .B1(new_n216), .B2(new_n218), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT73), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n219), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT76), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n209), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n223), .A2(new_n217), .B1(G101), .B2(new_n213), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n235), .A2(KEYINPUT5), .A3(G119), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n189), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT77), .A4(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT78), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n208), .B1(new_n229), .B2(new_n219), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n240), .B1(new_n247), .B2(new_n231), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n226), .A2(KEYINPUT76), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n244), .A2(KEYINPUT80), .A3(new_n245), .A4(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n250), .A2(new_n245), .A3(new_n243), .A4(new_n241), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT80), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n241), .A2(new_n243), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n226), .A2(KEYINPUT76), .B1(new_n233), .B2(new_n239), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT77), .B1(new_n258), .B2(new_n232), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n250), .A2(KEYINPUT79), .A3(new_n243), .A4(new_n241), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n248), .A2(new_n249), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n262), .B2(new_n242), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n265), .A2(KEYINPUT64), .A3(G146), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G128), .ZN(new_n273));
  INV_X1    g087(.A(new_n266), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n267), .ZN(new_n275));
  OAI21_X1  g089(.A(G128), .B1(new_n266), .B2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT0), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT0), .B(G128), .Z(new_n285));
  AOI22_X1  g099(.A1(new_n271), .A2(new_n284), .B1(new_n275), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G224), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT81), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n287), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n255), .A2(new_n264), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT84), .B1(new_n286), .B2(new_n280), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n287), .B(new_n295), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n213), .A2(G101), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n224), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT83), .B(new_n239), .C1(new_n298), .C2(KEYINPUT82), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n242), .B(KEYINPUT8), .Z(new_n300));
  OAI21_X1  g114(.A(KEYINPUT83), .B1(new_n298), .B2(KEYINPUT82), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n239), .B1(new_n233), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n262), .A2(new_n242), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n292), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n292), .A2(new_n307), .A3(new_n309), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT11), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G137), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT11), .A3(G134), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n316), .B(new_n318), .C1(G134), .C2(new_n317), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n319), .A2(G131), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n315), .A2(G137), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n317), .A2(G134), .ZN(new_n322));
  OAI21_X1  g136(.A(G131), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n278), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n319), .B(G131), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n286), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n327), .B2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n192), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n324), .A2(new_n191), .A3(new_n326), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n336));
  NOR2_X1   g150(.A1(G237), .A2(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G210), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G101), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n334), .A2(new_n335), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  INV_X1    g157(.A(new_n341), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n327), .A2(new_n192), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n335), .ZN(new_n347));
  INV_X1    g161(.A(new_n335), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT28), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n344), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n343), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G472), .ZN(new_n352));
  INV_X1    g166(.A(G902), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n335), .A4(new_n341), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n353), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n352), .A4(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n333), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n191), .B1(new_n362), .B2(new_n331), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(new_n348), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n341), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n347), .A2(new_n349), .A3(new_n344), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n353), .B1(new_n366), .B2(new_n367), .ZN(new_n370));
  OAI21_X1  g184(.A(G472), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n361), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  INV_X1    g187(.A(G140), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n280), .A2(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(G146), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G119), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G128), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(G128), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(KEYINPUT23), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(G110), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT24), .B(G110), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n385), .A2(KEYINPUT67), .A3(G128), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT67), .B1(new_n385), .B2(G128), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n386), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n384), .B(new_n393), .C1(new_n394), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n394), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n389), .B2(G110), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n378), .A2(G146), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n382), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT69), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT22), .B(G137), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n398), .B2(new_n403), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n353), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(KEYINPUT70), .A3(KEYINPUT25), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(G234), .B2(new_n353), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n409), .A2(new_n410), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n372), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n230), .A2(new_n286), .A3(new_n207), .ZN(new_n425));
  INV_X1    g239(.A(new_n325), .ZN(new_n426));
  INV_X1    g240(.A(new_n276), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n273), .B1(new_n271), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n233), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n278), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n425), .A2(new_n426), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n288), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n325), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n433), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n298), .A2(KEYINPUT74), .A3(new_n279), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n233), .B2(new_n278), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n446), .A3(new_n429), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n447), .B2(new_n325), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n325), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(KEYINPUT75), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n325), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n443), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n442), .B(G469), .C1(new_n454), .C2(new_n437), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n438), .B1(new_n450), .B2(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n437), .B1(new_n441), .B2(new_n433), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n456), .B(new_n353), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(new_n353), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT9), .B(G234), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n337), .A2(G214), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n265), .ZN(new_n467));
  AOI21_X1  g281(.A(G143), .B1(new_n337), .B2(G214), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G131), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n467), .A2(G131), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT17), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n382), .B(new_n383), .C1(new_n471), .C2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G113), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(new_n201), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(KEYINPUT90), .Z(new_n480));
  AOI21_X1  g294(.A(KEYINPUT85), .B1(new_n376), .B2(new_n377), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(G146), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n402), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n484), .B2(new_n402), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n469), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n469), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n486), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n492), .A2(new_n493), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT87), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n477), .B(new_n480), .C1(new_n495), .C2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n474), .A2(new_n476), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(KEYINPUT87), .A3(new_n498), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(new_n479), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n353), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G475), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n482), .A2(KEYINPUT19), .A3(new_n483), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n376), .A3(new_n377), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n510), .A3(new_n380), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT89), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n381), .B1(new_n471), .B2(new_n472), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n502), .A2(new_n503), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n500), .B1(new_n514), .B2(new_n479), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NOR2_X1   g330(.A1(G475), .A2(G902), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n507), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n521), .A2(G952), .A3(new_n288), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n235), .A2(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n527));
  INV_X1    g341(.A(G122), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G116), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n531));
  OAI21_X1  g345(.A(G107), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(G128), .B(G143), .Z(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(G134), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(G134), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n526), .A2(new_n529), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n536), .A2(new_n537), .B1(new_n198), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n198), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n538), .B(G107), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G128), .A3(new_n265), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(G134), .C1(new_n535), .C2(new_n546), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n545), .A3(new_n536), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  OR3_X1    g364(.A1(new_n463), .A2(new_n416), .A3(G953), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n353), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n555), .B(new_n557), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n520), .A2(new_n525), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n465), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n313), .A2(new_n423), .A3(new_n424), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G101), .ZN(G3));
  AND3_X1   g376(.A1(new_n292), .A2(new_n307), .A3(new_n309), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n309), .B1(new_n292), .B2(new_n307), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n424), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT94), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(new_n424), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n525), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n342), .A2(new_n343), .A3(new_n350), .ZN(new_n570));
  OAI21_X1  g384(.A(G472), .B1(new_n570), .B2(new_n357), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n571), .A2(new_n355), .ZN(new_n572));
  INV_X1    g386(.A(new_n422), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n465), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT33), .B1(new_n553), .B2(new_n554), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n550), .A2(new_n551), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n552), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n556), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n556), .A2(new_n353), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n555), .B2(G478), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n520), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n569), .A2(new_n575), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  OAI211_X1 g405(.A(new_n558), .B(new_n507), .C1(new_n518), .C2(new_n519), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n569), .A2(new_n575), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G107), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G9));
  NAND2_X1  g410(.A1(new_n398), .A2(new_n403), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n398), .A2(new_n599), .A3(new_n403), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(KEYINPUT36), .B2(new_n407), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n407), .A2(KEYINPUT36), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n598), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT97), .B1(new_n605), .B2(new_n421), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n602), .A2(new_n607), .A3(new_n420), .A4(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n418), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n571), .A2(new_n355), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n313), .A2(new_n560), .A3(new_n424), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT37), .B(G110), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  NAND2_X1  g429(.A1(new_n566), .A2(new_n568), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n610), .B1(new_n361), .B2(new_n371), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n465), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n522), .B1(new_n523), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n592), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n313), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n311), .A2(KEYINPUT38), .A3(new_n312), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n341), .B1(new_n346), .B2(new_n335), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT98), .Z(new_n631));
  INV_X1    g445(.A(new_n342), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n353), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n361), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n520), .A2(new_n558), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n636), .A2(new_n424), .A3(new_n610), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n622), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n462), .A2(new_n464), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT101), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n629), .B(new_n639), .C1(KEYINPUT40), .C2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(KEYINPUT40), .B2(new_n644), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G143), .ZN(G45));
  NOR2_X1   g461(.A1(new_n586), .A2(new_n622), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n620), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  OR2_X1    g464(.A1(new_n457), .A2(new_n458), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(G469), .B1(new_n652), .B2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n464), .A3(new_n459), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n654), .A2(new_n372), .A3(new_n422), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n569), .A2(new_n587), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G15));
  INV_X1    g472(.A(new_n525), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n616), .A2(new_n659), .A3(new_n593), .A4(new_n655), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  INV_X1    g475(.A(new_n654), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n618), .A2(new_n559), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n567), .B1(new_n313), .B2(new_n424), .ZN(new_n664));
  INV_X1    g478(.A(new_n568), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G119), .ZN(G21));
  NOR3_X1   g481(.A1(new_n654), .A2(new_n574), .A3(new_n525), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n638), .B(new_n668), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT102), .B(G122), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G24));
  AND2_X1   g485(.A1(new_n612), .A2(new_n648), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n616), .A2(new_n662), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G125), .ZN(G27));
  INV_X1    g488(.A(new_n424), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n563), .A2(new_n564), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n462), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n455), .A2(new_n459), .A3(KEYINPUT103), .A4(new_n461), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n678), .A2(new_n464), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n676), .A2(new_n680), .A3(new_n423), .A4(new_n648), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n311), .A2(new_n424), .A3(new_n312), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n678), .A2(new_n464), .A3(new_n679), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n423), .A4(new_n648), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n423), .B(KEYINPUT105), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(KEYINPUT42), .A3(new_n648), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G131), .ZN(G33));
  XNOR2_X1  g507(.A(new_n623), .B(KEYINPUT106), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n676), .A2(new_n680), .A3(new_n423), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G134), .ZN(G36));
  INV_X1    g510(.A(new_n459), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n450), .A2(new_n453), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n433), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(new_n436), .B1(new_n441), .B2(new_n439), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(KEYINPUT45), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n704), .A2(KEYINPUT108), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n461), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n697), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n461), .C1(new_n706), .C2(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n611), .A2(new_n609), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT111), .Z(new_n714));
  OR2_X1    g528(.A1(new_n581), .A2(new_n584), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n520), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n716), .B2(new_n520), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n585), .A2(KEYINPUT109), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n585), .A2(KEYINPUT109), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT43), .ZN(new_n721));
  INV_X1    g535(.A(new_n520), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n718), .A2(KEYINPUT43), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT44), .Z(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n684), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n712), .A2(new_n726), .A3(new_n464), .A4(new_n641), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G137), .ZN(G39));
  NAND2_X1  g542(.A1(new_n712), .A2(new_n464), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n372), .A2(new_n676), .A3(new_n422), .A4(new_n648), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  NAND2_X1  g550(.A1(new_n653), .A2(new_n459), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT49), .ZN(new_n738));
  INV_X1    g552(.A(new_n464), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n718), .A2(new_n675), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n636), .A2(new_n422), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n741), .B(new_n742), .C1(KEYINPUT49), .C2(new_n737), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n629), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n676), .A2(new_n662), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n718), .A2(KEYINPUT43), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n721), .A2(new_n722), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n522), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n723), .A2(KEYINPUT116), .A3(new_n522), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n690), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT48), .ZN(new_n757));
  INV_X1    g571(.A(new_n522), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n742), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n587), .ZN(new_n761));
  INV_X1    g575(.A(G952), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n574), .B1(new_n752), .B2(new_n753), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n654), .B1(new_n566), .B2(new_n568), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n762), .B(G953), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n757), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n756), .A2(KEYINPUT48), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n654), .A2(new_n424), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n629), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n771), .A2(KEYINPUT118), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n771), .B2(KEYINPUT118), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n722), .A2(new_n715), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n760), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n755), .A2(new_n612), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n769), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n760), .A2(new_n777), .B1(new_n755), .B2(new_n612), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(KEYINPUT120), .C1(new_n774), .C2(new_n773), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n763), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n684), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT47), .B1(new_n712), .B2(new_n464), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n730), .B(new_n739), .C1(new_n710), .C2(new_n711), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n737), .A2(new_n464), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n768), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n656), .A2(new_n660), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n525), .B1(new_n586), .B2(new_n592), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n313), .A2(new_n424), .A3(new_n575), .A4(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n561), .A2(new_n613), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n666), .A3(new_n669), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  OAI221_X1 g615(.A(new_n619), .B1(new_n623), .B2(new_n648), .C1(new_n664), .C2(new_n665), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n609), .A2(new_n622), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT113), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n680), .A2(new_n635), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n616), .A2(new_n638), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n673), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n686), .A2(new_n672), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n520), .A2(new_n558), .A3(new_n622), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n617), .A2(new_n464), .A3(new_n462), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n812), .B2(new_n676), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n684), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n809), .B(new_n695), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n689), .B2(new_n691), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n802), .A2(new_n673), .A3(new_n806), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n801), .A2(new_n808), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n795), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n808), .A2(new_n819), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n799), .A2(new_n666), .A3(new_n669), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n569), .B(new_n655), .C1(new_n587), .C2(new_n593), .ZN(new_n825));
  INV_X1    g639(.A(new_n816), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n692), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n827), .A3(KEYINPUT114), .A4(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n821), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n827), .A3(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n829), .A3(KEYINPUT115), .A4(new_n833), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n787), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT117), .B(new_n786), .C1(new_n733), .C2(new_n791), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n775), .A2(new_n780), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n794), .B(new_n838), .C1(new_n839), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(G952), .A2(G953), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n744), .B1(new_n846), .B2(new_n847), .ZN(G75));
  NOR2_X1   g662(.A1(new_n288), .A2(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n353), .B1(new_n832), .B2(new_n829), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT56), .B1(new_n851), .B2(G210), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n255), .A2(new_n264), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n291), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT55), .Z(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n852), .B2(new_n855), .ZN(G51));
  NAND2_X1  g671(.A1(new_n832), .A2(new_n829), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n834), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n460), .B(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n652), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n706), .A2(new_n707), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n851), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n849), .B1(new_n865), .B2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  INV_X1    g683(.A(new_n515), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n849), .ZN(G60));
  XOR2_X1   g687(.A(new_n582), .B(KEYINPUT59), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n838), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n580), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(KEYINPUT123), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n580), .A2(new_n874), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n859), .B2(new_n834), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT122), .B1(new_n879), .B2(new_n849), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n832), .A2(new_n829), .A3(new_n833), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n833), .B1(new_n832), .B2(new_n829), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n881), .B(new_n850), .C1(new_n884), .C2(new_n878), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT123), .B1(new_n875), .B2(new_n876), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(G63));
  NAND2_X1  g703(.A1(G217), .A2(G902), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT60), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n858), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n849), .B1(new_n892), .B2(new_n419), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n605), .B2(new_n892), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g709(.A1(G224), .A2(G953), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n524), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n801), .B2(new_n288), .ZN(new_n898));
  INV_X1    g712(.A(G898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n853), .B1(new_n899), .B2(G953), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n898), .B(new_n900), .Z(G69));
  AND3_X1   g715(.A1(new_n616), .A2(new_n690), .A3(new_n638), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n712), .A2(new_n464), .A3(new_n641), .A4(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n802), .A2(new_n673), .A3(new_n695), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n727), .A2(new_n692), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n735), .A2(new_n288), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n362), .A2(new_n331), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n508), .A2(new_n510), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(new_n910));
  OAI211_X1 g724(.A(new_n906), .B(new_n910), .C1(new_n621), .C2(new_n288), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n646), .A2(new_n673), .A3(new_n802), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n586), .A2(new_n592), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT125), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n643), .A2(new_n423), .A3(new_n676), .A4(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n727), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n735), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n288), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n911), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G72));
  NOR2_X1   g737(.A1(new_n364), .A2(new_n344), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n914), .A2(new_n735), .A3(new_n801), .A4(new_n918), .ZN(new_n926));
  NAND2_X1  g740(.A1(G472), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT63), .Z(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT126), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n632), .A2(KEYINPUT127), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n365), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n830), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n928), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n735), .A2(new_n903), .A3(new_n905), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n801), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n364), .A2(new_n344), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n933), .B(new_n850), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n930), .A2(new_n938), .ZN(G57));
endmodule


