//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(new_n194), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n189), .A3(new_n197), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n190), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n188), .B2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n202), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G224), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n214), .A2(new_n216), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(G104), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n222), .A2(new_n228), .A3(new_n223), .A4(G104), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT77), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n230), .A2(G101), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(G101), .ZN(new_n234));
  INV_X1    g048(.A(G101), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n225), .A2(new_n235), .A3(new_n227), .A4(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n232), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n244), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT83), .B1(new_n238), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(G110), .B(G122), .Z(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n246), .ZN(new_n251));
  INV_X1    g065(.A(G113), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n253));
  INV_X1    g067(.A(new_n240), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n253), .A2(new_n243), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n223), .A2(G104), .ZN(new_n259));
  OAI21_X1  g073(.A(G101), .B1(new_n259), .B2(new_n226), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n236), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n237), .A2(new_n234), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n230), .A2(G101), .A3(new_n232), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  INV_X1    g080(.A(new_n247), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n248), .A2(new_n250), .A3(new_n262), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n272));
  AOI211_X1 g086(.A(KEYINPUT83), .B(new_n247), .C1(new_n263), .C2(new_n264), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT85), .A3(new_n250), .A4(new_n262), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n262), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n249), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n221), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(new_n277), .B2(new_n249), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n220), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n214), .B1(KEYINPUT7), .B2(new_n216), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n271), .B2(new_n275), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n249), .A2(KEYINPUT8), .ZN(new_n285));
  INV_X1    g099(.A(new_n261), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n258), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT5), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n251), .B1(new_n256), .B2(new_n288), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n285), .B(new_n287), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n249), .A2(KEYINPUT8), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n290), .A2(new_n291), .B1(KEYINPUT7), .B2(new_n217), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n281), .A2(new_n282), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n282), .B1(new_n281), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT86), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n298), .B(new_n187), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n203), .A2(new_n189), .A3(new_n197), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G128), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n193), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n261), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n200), .B2(new_n265), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n311));
  INV_X1    g125(.A(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G134), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT65), .A3(G137), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT11), .B1(new_n312), .B2(G134), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(G137), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G131), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n316), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n312), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n325), .B2(new_n316), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n305), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n189), .A2(KEYINPUT78), .A3(KEYINPUT1), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(G128), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n304), .B1(new_n332), .B2(new_n198), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n308), .B1(new_n333), .B2(new_n261), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n310), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G140), .ZN(new_n336));
  INV_X1    g150(.A(G227), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G953), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n336), .B(new_n338), .Z(new_n339));
  AND2_X1   g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n310), .A2(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n327), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n333), .A2(new_n261), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n211), .B1(new_n236), .B2(new_n260), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT12), .B(new_n327), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT79), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n327), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT12), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n261), .A2(new_n307), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n261), .B2(new_n333), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT12), .A4(new_n327), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n348), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(new_n335), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n356), .B2(new_n335), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n339), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n344), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n303), .B1(new_n362), .B2(G469), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(KEYINPUT81), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n348), .A2(new_n351), .A3(new_n365), .A4(new_n355), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n340), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT82), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n335), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n361), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n364), .A2(new_n340), .A3(new_n371), .A4(new_n366), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n301), .A3(new_n302), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n239), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n202), .A2(G119), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT24), .B(G110), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n384), .B2(G110), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n386));
  XNOR2_X1  g200(.A(G125), .B(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n188), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n188), .B(new_n389), .C1(KEYINPUT16), .C2(new_n387), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(new_n380), .C1(new_n384), .C2(G110), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n386), .A2(new_n388), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n384), .A2(G110), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n396));
  INV_X1    g210(.A(new_n389), .ZN(new_n397));
  AOI21_X1  g211(.A(G146), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI221_X1 g212(.A(new_n395), .B1(new_n378), .B2(new_n379), .C1(new_n390), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT22), .B(G137), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n399), .A3(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(G234), .B2(new_n302), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(G902), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT75), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n405), .A2(new_n302), .A3(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT73), .B1(new_n414), .B2(KEYINPUT25), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT25), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT74), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n420), .A3(new_n418), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n417), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n412), .B1(new_n422), .B2(new_n409), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT9), .B(G234), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n425), .B2(G902), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n375), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n199), .B(new_n196), .C1(new_n323), .C2(new_n326), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n312), .A2(G134), .ZN(new_n431));
  OAI21_X1  g245(.A(G131), .B1(new_n319), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n211), .A2(new_n322), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n434), .B2(new_n267), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n267), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n322), .A2(new_n432), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT66), .B1(new_n437), .B2(new_n307), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT66), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n211), .A2(new_n439), .A3(new_n322), .A4(new_n432), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n430), .A3(new_n247), .A4(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n435), .B(new_n436), .C1(new_n429), .C2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G237), .A2(G953), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G210), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(G101), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n430), .A2(new_n450), .A3(new_n433), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n438), .A2(new_n430), .A3(new_n440), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(KEYINPUT30), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n447), .B(new_n441), .C1(new_n453), .C2(new_n247), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n454), .B2(KEYINPUT31), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n430), .A2(new_n450), .A3(new_n433), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n247), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n441), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n458), .A2(new_n448), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT67), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n463), .A3(KEYINPUT31), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n455), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G472), .A2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n428), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n267), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT70), .A3(new_n441), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n452), .A2(new_n471), .A3(new_n267), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(KEYINPUT28), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT29), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n448), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n435), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n476), .A2(new_n302), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n459), .A2(KEYINPUT28), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n447), .A3(new_n436), .A4(new_n435), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n456), .A2(new_n457), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n459), .B1(new_n480), .B2(new_n267), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n474), .B(new_n479), .C1(new_n481), .C2(new_n447), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n485), .A2(KEYINPUT69), .A3(new_n474), .A4(new_n479), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n477), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G472), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n460), .A2(new_n461), .B1(new_n448), .B2(new_n442), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n454), .A2(new_n463), .A3(KEYINPUT31), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n463), .B1(new_n454), .B2(KEYINPUT31), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT32), .A3(new_n466), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n468), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT71), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n468), .A2(new_n488), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n427), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n390), .A2(new_n398), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n443), .A2(G143), .A3(G214), .ZN(new_n500));
  AOI21_X1  g314(.A(G143), .B1(new_n443), .B2(G214), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT17), .B(G131), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT89), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n500), .A2(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n321), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n500), .B2(new_n501), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n499), .B(new_n514), .C1(new_n504), .C2(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n507), .A2(new_n513), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n508), .B1(new_n518), .B2(new_n321), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n387), .B(new_n188), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(new_n518), .C2(new_n510), .ZN(new_n521));
  XNOR2_X1  g335(.A(G113), .B(G122), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT87), .B(G104), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n387), .B(KEYINPUT19), .Z(new_n527));
  OAI21_X1  g341(.A(new_n391), .B1(new_n527), .B2(G146), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n509), .A2(new_n510), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n524), .ZN(new_n531));
  AOI21_X1  g345(.A(G475), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT91), .B1(new_n526), .B2(new_n531), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT20), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n302), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n525), .B1(new_n517), .B2(new_n521), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n302), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G475), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n532), .A2(new_n534), .A3(new_n302), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n532), .B2(new_n302), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n526), .A2(new_n531), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n544), .B(new_n545), .C1(G475), .C2(G902), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(G234), .A2(G237), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(G952), .A3(new_n215), .ZN(new_n549));
  XOR2_X1   g363(.A(KEYINPUT21), .B(G898), .Z(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(G902), .A3(G953), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n241), .A2(G122), .ZN(new_n553));
  INV_X1    g367(.A(G122), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT92), .B1(new_n554), .B2(G116), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n241), .A3(G122), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n223), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(new_n553), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n190), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n202), .A2(G143), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n314), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n558), .B1(KEYINPUT14), .B2(new_n223), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n569), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n190), .A2(KEYINPUT93), .A3(KEYINPUT13), .A4(G128), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(new_n563), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G134), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n564), .A2(new_n314), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n558), .A2(new_n223), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n575), .C1(new_n559), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n425), .A2(new_n408), .A3(G953), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT94), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n582), .B(new_n584), .Z(new_n585));
  NAND3_X1  g399(.A1(new_n547), .A2(new_n552), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n300), .A2(new_n498), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(new_n426), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n363), .B2(new_n374), .ZN(new_n591));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n492), .B2(new_n302), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n465), .A2(new_n467), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n423), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n187), .B(new_n552), .C1(new_n294), .C2(new_n295), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n580), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n580), .A2(new_n598), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(G478), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(G478), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n581), .A2(new_n583), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NOR4_X1   g418(.A1(new_n596), .A2(new_n597), .A3(new_n547), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT34), .B(G104), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  AOI21_X1  g421(.A(new_n543), .B1(G475), .B2(new_n538), .ZN(new_n608));
  INV_X1    g422(.A(new_n585), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n596), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT35), .B(G107), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NAND2_X1  g427(.A1(new_n422), .A2(new_n409), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n404), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n400), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n617), .A2(new_n411), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n375), .A2(new_n426), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n300), .A2(new_n587), .A3(new_n595), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G110), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  NOR2_X1   g439(.A1(new_n620), .A2(new_n296), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n495), .A2(new_n497), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n551), .A2(G900), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n549), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n610), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT96), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n626), .A2(new_n627), .A3(new_n634), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  NOR2_X1   g451(.A1(new_n294), .A2(new_n295), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT38), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n281), .A2(new_n293), .ZN(new_n640));
  INV_X1    g454(.A(new_n282), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n281), .A2(new_n282), .A3(new_n293), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n187), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n532), .A2(new_n302), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT20), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n532), .A2(new_n534), .A3(new_n302), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n546), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n535), .A2(new_n539), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n609), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n481), .A2(new_n448), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n447), .B1(new_n470), .B2(new_n472), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n302), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n657), .A2(new_n656), .A3(new_n658), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n468), .A3(new_n493), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n647), .A2(new_n648), .A3(new_n655), .A4(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n619), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n629), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n591), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n666), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  INV_X1    g486(.A(new_n604), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n654), .A2(new_n673), .A3(new_n629), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n626), .A2(new_n627), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT98), .B(G146), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G48));
  INV_X1    g492(.A(new_n423), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n495), .B2(new_n497), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n547), .A2(new_n604), .ZN(new_n681));
  INV_X1    g495(.A(new_n597), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n373), .A2(new_n302), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n426), .A3(new_n374), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n680), .A2(new_n681), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NOR2_X1   g503(.A1(new_n597), .A2(new_n610), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n690), .A3(new_n686), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  AOI21_X1  g506(.A(new_n586), .B1(new_n495), .B2(new_n497), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n296), .A2(new_n685), .A3(new_n666), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT99), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NOR2_X1   g514(.A1(new_n655), .A2(KEYINPUT102), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n654), .B2(new_n609), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n593), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  INV_X1    g520(.A(new_n412), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n614), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g522(.A(KEYINPUT101), .B(new_n412), .C1(new_n422), .C2(new_n409), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n460), .A2(new_n461), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n454), .A2(KEYINPUT31), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n473), .A2(new_n435), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n447), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n466), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n705), .A2(new_n710), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n704), .A2(new_n718), .A3(new_n682), .A4(new_n686), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(G122), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G24));
  NOR2_X1   g535(.A1(new_n296), .A2(new_n685), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n705), .A2(new_n717), .A3(new_n619), .A4(new_n716), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n675), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(new_n591), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n642), .A2(new_n187), .A3(new_n643), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n726), .A2(new_n727), .A3(new_n674), .ZN(new_n728));
  INV_X1    g542(.A(new_n710), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n488), .A2(new_n493), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(new_n732), .A3(KEYINPUT42), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT42), .B1(new_n728), .B2(new_n680), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g550(.A(KEYINPUT104), .B(KEYINPUT42), .C1(new_n728), .C2(new_n680), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(new_n727), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n498), .A2(new_n631), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(new_n595), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n547), .B2(new_n673), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n652), .A2(new_n653), .A3(new_n673), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n743), .B(new_n619), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n747), .B1(KEYINPUT107), .B2(new_n744), .ZN(new_n753));
  INV_X1    g567(.A(new_n748), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n547), .A2(new_n673), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n595), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n619), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n752), .A2(new_n757), .A3(new_n740), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n356), .A2(new_n335), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT80), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n356), .A2(new_n357), .A3(new_n335), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n361), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT45), .A3(new_n343), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT105), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n765), .A3(KEYINPUT45), .A4(new_n343), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n362), .A2(KEYINPUT45), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n303), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n303), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n769), .A2(KEYINPUT106), .A3(KEYINPUT46), .A4(new_n770), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n776), .A3(new_n374), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n758), .A2(new_n426), .A3(new_n667), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NOR4_X1   g594(.A1(new_n627), .A2(new_n423), .A3(new_n674), .A4(new_n727), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n426), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT47), .B1(new_n778), .B2(new_n426), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n676), .A2(new_n724), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n635), .B2(new_n633), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n701), .A2(new_n296), .A3(new_n703), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n619), .A2(new_n630), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n591), .A3(new_n663), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n790), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n791), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n790), .A2(new_n636), .A3(new_n797), .A4(new_n795), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n687), .A2(new_n719), .A3(new_n691), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n552), .A2(new_n591), .A3(new_n595), .A4(new_n423), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n300), .A2(new_n681), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n588), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n588), .B2(new_n802), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n800), .B(new_n699), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n654), .A2(new_n585), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n300), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n622), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(new_n622), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n620), .A2(new_n609), .A3(new_n630), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n627), .A3(new_n608), .A4(new_n740), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n728), .A2(new_n723), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n738), .A2(new_n741), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n799), .A2(KEYINPUT53), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n813), .A2(new_n818), .ZN(new_n822));
  INV_X1    g636(.A(new_n796), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n792), .A2(new_n790), .A3(new_n795), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n811), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n809), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n687), .A2(new_n719), .A3(new_n691), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n698), .B2(new_n696), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n588), .A2(new_n802), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n588), .A2(new_n802), .A3(new_n803), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n738), .A2(new_n741), .A3(new_n817), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT53), .A4(new_n799), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n826), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n842), .A3(new_n819), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n549), .B1(new_n753), .B2(new_n755), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n718), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n187), .B1(new_n639), .B2(new_n646), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(KEYINPUT50), .A3(new_n686), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n718), .A2(new_n844), .A3(new_n686), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n647), .A2(new_n648), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n847), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n663), .A2(new_n549), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n740), .A2(new_n854), .A3(new_n686), .A4(new_n423), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n654), .A3(new_n673), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n844), .A2(new_n686), .A3(new_n740), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n723), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n852), .B1(new_n847), .B2(new_n851), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n778), .A2(new_n426), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT47), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n426), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n684), .A2(new_n374), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n590), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n740), .A3(new_n845), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT51), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n845), .A2(new_n722), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n732), .A2(new_n844), .A3(new_n686), .A4(new_n740), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT48), .A3(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n855), .A2(new_n547), .A3(new_n604), .ZN(new_n876));
  INV_X1    g690(.A(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(G953), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n875), .B(new_n878), .C1(KEYINPUT48), .C2(new_n874), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n847), .A2(new_n851), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n858), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n869), .A2(KEYINPUT51), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n869), .A2(KEYINPUT114), .A3(KEYINPUT51), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n841), .A2(new_n843), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n877), .A2(new_n215), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n841), .A2(new_n888), .A3(new_n892), .A4(new_n843), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n729), .A2(new_n648), .A3(new_n590), .A4(new_n747), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT109), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n866), .B(KEYINPUT49), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n647), .A3(new_n664), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n302), .B1(new_n826), .B2(new_n819), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n279), .A2(new_n280), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n220), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n215), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n900), .A2(new_n775), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT117), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n303), .B(KEYINPUT57), .ZN(new_n912));
  INV_X1    g726(.A(new_n843), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n842), .B1(new_n826), .B2(new_n819), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n373), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n908), .B1(new_n911), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n918), .A2(new_n526), .A3(new_n531), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n526), .B2(new_n531), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n908), .ZN(G60));
  INV_X1    g735(.A(new_n908), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n599), .A2(new_n600), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n602), .B(KEYINPUT59), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n923), .B(new_n925), .C1(new_n913), .C2(new_n914), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n841), .B2(new_n843), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n922), .B(new_n926), .C1(new_n927), .C2(new_n923), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(G63));
  NOR2_X1   g743(.A1(new_n408), .A2(new_n302), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n932), .B(new_n934), .C1(new_n826), .C2(new_n819), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n908), .B1(new_n935), .B2(new_n616), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n939));
  INV_X1    g753(.A(new_n932), .ZN(new_n940));
  INV_X1    g754(.A(new_n819), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n837), .B2(new_n799), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n940), .B(new_n933), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n407), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n922), .B1(new_n943), .B2(new_n617), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n934), .B1(new_n826), .B2(new_n819), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n947), .A2(new_n940), .B1(new_n406), .B2(new_n405), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n937), .B(KEYINPUT61), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n945), .A2(new_n949), .ZN(G66));
  AOI21_X1  g764(.A(new_n215), .B1(new_n550), .B2(G224), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT119), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n835), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n828), .A2(new_n830), .A3(new_n834), .A4(KEYINPUT119), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n955), .B2(new_n215), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n903), .B1(G898), .B2(new_n215), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  INV_X1    g772(.A(G900), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n337), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT121), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n793), .A2(new_n732), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(new_n426), .A3(new_n667), .A4(new_n778), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n779), .A2(new_n792), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n738), .A2(new_n741), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n788), .A2(new_n966), .A3(new_n215), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n453), .B(KEYINPUT120), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n527), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n792), .A2(new_n671), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n681), .A2(new_n807), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(new_n668), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n680), .A3(new_n740), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n977), .A2(new_n779), .A3(new_n788), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n969), .B1(new_n981), .B2(new_n215), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n961), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n961), .B(KEYINPUT122), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n972), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT124), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n961), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n972), .B(KEYINPUT123), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n982), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n992), .A3(new_n986), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n481), .A2(new_n448), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n657), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n840), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n996), .B(KEYINPUT125), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n981), .B2(new_n955), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n657), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n953), .A2(new_n788), .A3(new_n966), .A4(new_n954), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n997), .B1(new_n1006), .B2(new_n1002), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT126), .B1(new_n1007), .B2(new_n908), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1007), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n922), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(new_n1000), .A3(new_n1008), .A4(new_n1004), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(G57));
endmodule


