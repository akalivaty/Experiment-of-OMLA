//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  NOR4_X1   g0024(.A1(new_n217), .A2(new_n220), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n209), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g0036(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G20), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(G1), .A2(G13), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(G50), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  AOI211_X1 g0043(.A(new_n212), .B(new_n235), .C1(new_n241), .C2(new_n243), .ZN(G361));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n227), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT2), .B(G226), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G264), .B(G270), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G358));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(G87), .B(G97), .Z(new_n256));
  XNOR2_X1  g0056(.A(G107), .B(G116), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n255), .B(new_n258), .ZN(G351));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G223), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT66), .B(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n260), .B1(new_n261), .B2(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n265), .B(new_n269), .C1(G77), .C2(new_n260), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n271), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n270), .B(new_n273), .C1(new_n219), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G179), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT69), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G58), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n239), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n289));
  OAI221_X1 g0089(.A(KEYINPUT68), .B1(new_n283), .B2(new_n285), .C1(new_n281), .C2(new_n282), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n240), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n291), .A2(new_n293), .B1(new_n218), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n206), .B2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G50), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n275), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n277), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n296), .A2(KEYINPUT9), .A3(new_n298), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n275), .A2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n275), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n305), .A2(new_n309), .A3(new_n306), .A4(new_n311), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n303), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n260), .B1(new_n232), .B2(new_n262), .C1(new_n263), .C2(new_n227), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT70), .B(G107), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n269), .C1(new_n318), .C2(new_n260), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n273), .C1(new_n214), .C2(new_n274), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n320), .B(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT8), .B(G58), .Z(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT65), .B(G20), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n284), .B1(new_n325), .B2(G77), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n282), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n293), .B1(new_n213), .B2(new_n295), .ZN(new_n330));
  INV_X1    g0130(.A(new_n297), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n213), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n323), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n322), .B2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n322), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n315), .A2(new_n316), .A3(new_n336), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n274), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G238), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n266), .A2(new_n215), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G232), .A2(G1698), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n263), .B2(new_n219), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n260), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n273), .B(new_n342), .C1(new_n346), .C2(new_n268), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G33), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT66), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G226), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n352), .B1(new_n357), .B2(new_n344), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n269), .B1(new_n358), .B2(new_n343), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n273), .A4(new_n342), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n348), .A2(new_n361), .A3(KEYINPUT73), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n347), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(G169), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(KEYINPUT14), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n348), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n348), .B1(new_n367), .B2(new_n361), .ZN(new_n370));
  OAI21_X1  g0170(.A(G179), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n362), .A2(new_n363), .A3(G169), .A4(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n366), .A2(new_n371), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT12), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n295), .B2(new_n231), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n294), .A2(KEYINPUT12), .A3(G68), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n331), .A2(new_n231), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n284), .A2(G50), .ZN(new_n380));
  XOR2_X1   g0180(.A(new_n380), .B(KEYINPUT75), .Z(new_n381));
  OAI221_X1 g0181(.A(new_n381), .B1(new_n207), .B2(G68), .C1(new_n213), .C2(new_n282), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n293), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n385), .A3(new_n293), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n379), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n375), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n362), .A2(new_n363), .A3(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n361), .A2(new_n367), .ZN(new_n393));
  INV_X1    g0193(.A(new_n348), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n310), .B1(new_n395), .B2(new_n368), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n390), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G190), .B1(new_n369), .B2(new_n370), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n391), .A4(new_n387), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n389), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n340), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n293), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n260), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n239), .A2(new_n352), .A3(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G68), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n226), .A2(new_n231), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n410), .B2(new_n202), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n284), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n404), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n239), .A2(new_n405), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n266), .A3(KEYINPUT3), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT78), .B1(new_n350), .B2(G33), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n350), .A2(G33), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n420), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n421), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n349), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n420), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n419), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n405), .B1(new_n431), .B2(new_n207), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(G68), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n417), .A2(new_n435), .ZN(new_n436));
  MUX2_X1   g0236(.A(new_n331), .B(new_n294), .S(new_n281), .Z(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n341), .A2(G232), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n263), .A2(new_n261), .B1(new_n219), .B2(new_n262), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n350), .A2(KEYINPUT78), .A3(G33), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n349), .B2(new_n427), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n440), .A2(new_n442), .B1(G33), .B2(G87), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n439), .B(new_n273), .C1(new_n443), .C2(new_n268), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n444), .A2(new_n334), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(G169), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n448), .B(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n444), .A2(new_n310), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n436), .A2(new_n451), .A3(new_n437), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n315), .A2(new_n336), .A3(new_n339), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT72), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n403), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n206), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n404), .A2(new_n294), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n327), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n237), .A2(G20), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n466));
  OAI211_X1 g0266(.A(G33), .B(G97), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n266), .A3(new_n215), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n221), .A2(new_n215), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n325), .B1(new_n318), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n428), .A2(G68), .A3(new_n239), .A4(new_n422), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n293), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n327), .A2(new_n294), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n464), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g0278(.A(KEYINPUT81), .B(new_n476), .C1(new_n474), .C2(new_n293), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n463), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n268), .B(G250), .C1(G1), .C2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n483), .A2(new_n272), .A3(G1), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n263), .A2(new_n232), .B1(new_n214), .B2(new_n262), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n442), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n484), .B(new_n486), .C1(new_n490), .C2(new_n268), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G169), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n334), .B2(new_n491), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT82), .B(new_n463), .C1(new_n478), .C2(new_n479), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n478), .A2(new_n479), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(G200), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n462), .A2(G87), .ZN(new_n498));
  INV_X1    g0298(.A(new_n491), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G190), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT83), .B1(new_n495), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n221), .B1(new_n236), .B2(new_n238), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n260), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n236), .A2(new_n238), .A3(new_n228), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n228), .A2(KEYINPUT70), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n228), .A2(KEYINPUT70), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT23), .B(G20), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n488), .A2(new_n207), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n505), .A2(new_n428), .A3(KEYINPUT22), .A4(new_n422), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n508), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n506), .A2(new_n507), .B1(new_n207), .B2(new_n488), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n515), .A4(new_n517), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n293), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n462), .A2(G107), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n294), .A2(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT25), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT5), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n206), .B(G45), .C1(new_n529), .C2(G41), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n530), .A2(new_n272), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n268), .B(G264), .C1(new_n530), .C2(new_n531), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n263), .A2(new_n222), .B1(new_n216), .B2(new_n262), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n442), .B1(G33), .B2(G294), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n533), .B(new_n534), .C1(new_n536), .C2(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G169), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  INV_X1    g0339(.A(new_n537), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G179), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(new_n542), .A3(G169), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n528), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n523), .A2(new_n293), .B1(G107), .B2(new_n462), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n535), .A2(new_n442), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n269), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n550), .A2(new_n310), .A3(new_n533), .A4(new_n534), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n537), .A2(new_n338), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT86), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT86), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n540), .A2(new_n554), .A3(new_n310), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n546), .A2(new_n527), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n545), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n268), .B(G270), .C1(new_n530), .C2(new_n531), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT84), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n229), .A2(new_n262), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n431), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n352), .A2(G303), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n428), .A2(G257), .A3(new_n422), .A4(new_n356), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n428), .A2(KEYINPUT84), .A3(new_n422), .A4(new_n561), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n567), .B2(new_n269), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G190), .A3(new_n533), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n462), .A2(G116), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n295), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G283), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n266), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n215), .A2(G33), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n325), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(G20), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n293), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n574), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n239), .C1(G33), .C2(new_n215), .ZN(new_n582));
  INV_X1    g0382(.A(new_n579), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT20), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n570), .B(new_n572), .C1(new_n580), .C2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI211_X1 g0386(.A(new_n559), .B(new_n532), .C1(new_n567), .C2(new_n269), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n569), .B(new_n586), .C1(new_n338), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(G179), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(G169), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n590), .A2(new_n587), .A3(KEYINPUT21), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n568), .A2(new_n533), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n571), .B2(new_n295), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n300), .B1(new_n596), .B2(new_n570), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n592), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n588), .B(new_n589), .C1(new_n591), .C2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n408), .A2(new_n318), .B1(G77), .B2(new_n284), .ZN(new_n600));
  XOR2_X1   g0400(.A(KEYINPUT80), .B(G107), .Z(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(KEYINPUT6), .B2(G97), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n601), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n325), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n293), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n462), .A2(G97), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n294), .A2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n268), .B1(new_n530), .B2(new_n531), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(new_n216), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n581), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT4), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n214), .B1(new_n353), .B2(new_n355), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n422), .A4(new_n428), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n260), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n269), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n300), .B1(new_n623), .B2(new_n533), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n260), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT4), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n619), .A2(new_n428), .A3(new_n618), .A4(new_n422), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n616), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n533), .B(new_n613), .C1(new_n628), .C2(new_n268), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n334), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n611), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(G190), .A3(new_n533), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(G200), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n609), .B1(new_n606), .B2(new_n293), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n608), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n557), .A2(new_n599), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n504), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n459), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT87), .Z(G372));
  INV_X1    g0440(.A(new_n336), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n400), .A2(new_n641), .B1(new_n388), .B2(new_n375), .ZN(new_n642));
  INV_X1    g0442(.A(new_n454), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n450), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n312), .A2(new_n314), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n303), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT89), .B1(new_n624), .B2(new_n630), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(G169), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n648), .B(new_n649), .C1(new_n334), .C2(new_n629), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n611), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT90), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n497), .A2(KEYINPUT88), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n491), .A2(new_n655), .A3(G200), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n496), .A3(new_n498), .A4(new_n500), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n480), .A2(new_n493), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n647), .A2(KEYINPUT90), .A3(new_n650), .A4(new_n611), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n653), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n589), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT21), .B1(new_n590), .B2(new_n587), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n593), .A2(new_n597), .A3(new_n592), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n545), .ZN(new_n668));
  INV_X1    g0468(.A(new_n636), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n556), .A3(new_n669), .A4(new_n658), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n663), .A2(new_n670), .A3(new_n659), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n495), .A2(new_n501), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT83), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n501), .ZN(new_n676));
  INV_X1    g0476(.A(new_n631), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n646), .B1(new_n459), .B2(new_n681), .ZN(G369));
  INV_X1    g0482(.A(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n325), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT27), .B1(new_n685), .B2(G1), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n687), .A3(new_n206), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n689), .A2(KEYINPUT91), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT91), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n586), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n589), .B1(new_n591), .B2(new_n598), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n599), .A2(new_n695), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n528), .A2(new_n693), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n557), .A2(new_n702), .B1(new_n545), .B2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n667), .B2(new_n693), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n694), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n545), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n703), .B1(new_n709), .B2(new_n694), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n210), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n318), .A2(G116), .A3(new_n471), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n713), .A2(new_n206), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT93), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  INV_X1    g0519(.A(new_n713), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n242), .C2(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n722));
  XNOR2_X1  g0522(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n629), .A2(new_n537), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n499), .B1(new_n724), .B2(KEYINPUT95), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n629), .A2(new_n726), .A3(new_n537), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n334), .A3(new_n593), .A4(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n622), .A2(new_n269), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n568), .A2(new_n731), .A3(new_n533), .A4(new_n613), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n540), .A2(new_n499), .A3(G179), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n537), .A2(new_n491), .A3(new_n334), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n587), .A4(new_n623), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n693), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n734), .A2(new_n736), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n728), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n693), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n637), .A2(new_n675), .A3(new_n676), .A4(new_n694), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n700), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT96), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(KEYINPUT96), .B(new_n700), .C1(new_n744), .C2(new_n745), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n675), .A2(new_n661), .A3(new_n676), .A4(new_n677), .ZN(new_n751));
  INV_X1    g0551(.A(new_n659), .ZN(new_n752));
  AND4_X1   g0552(.A1(new_n556), .A2(new_n658), .A3(new_n631), .A4(new_n635), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n668), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n653), .A2(new_n660), .A3(new_n662), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n751), .B(new_n754), .C1(new_n661), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n693), .B1(new_n672), .B2(new_n679), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(KEYINPUT29), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n750), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n723), .B1(new_n760), .B2(G1), .ZN(G364));
  OAI21_X1  g0561(.A(G1), .B1(new_n685), .B2(new_n483), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n713), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n701), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n699), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(G330), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n240), .B1(G20), .B2(new_n300), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n310), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n239), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n239), .A2(new_n334), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT97), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n775), .A3(G200), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n774), .A2(new_n310), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n771), .B1(new_n777), .B2(new_n231), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT99), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n338), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n325), .A2(new_n310), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n228), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n239), .A2(new_n334), .A3(G190), .A4(G200), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G77), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n774), .A2(G190), .A3(new_n776), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n779), .B(new_n784), .C1(new_n218), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n772), .A2(G190), .A3(new_n338), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n260), .B1(new_n787), .B2(new_n226), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n780), .A2(G20), .A3(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n221), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n239), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G159), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  INV_X1    g0597(.A(new_n783), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n785), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n777), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n787), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G322), .ZN(new_n804));
  INV_X1    g0604(.A(new_n781), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G329), .A2(new_n791), .B1(new_n805), .B2(G283), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n260), .B1(new_n770), .B2(G294), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n804), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n789), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n799), .B(new_n808), .C1(G303), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n767), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n431), .A2(KEYINPUT79), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n425), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n712), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n243), .A2(new_n483), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n483), .C2(new_n255), .ZN(new_n817));
  INV_X1    g0617(.A(G355), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n210), .A2(new_n260), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(G116), .B2(new_n210), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n767), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n811), .A2(new_n763), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT100), .Z(new_n827));
  INV_X1    g0627(.A(new_n823), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n765), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n766), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0631(.A1(new_n336), .A2(new_n693), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n339), .B1(new_n333), .B2(new_n694), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n336), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n758), .B(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n745), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n742), .B1(new_n741), .B2(new_n693), .ZN(new_n838));
  AOI211_X1 g0638(.A(KEYINPUT31), .B(new_n694), .C1(new_n740), .C2(new_n728), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(G330), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT96), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n746), .A2(new_n747), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n836), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT102), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n763), .B1(new_n836), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n352), .B1(new_n789), .B2(new_n228), .ZN(new_n849));
  INV_X1    g0649(.A(G294), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n787), .A2(new_n850), .B1(new_n221), .B2(new_n781), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G116), .C2(new_n783), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n800), .A2(G283), .B1(G311), .B2(new_n791), .ZN(new_n853));
  INV_X1    g0653(.A(new_n785), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G303), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(new_n771), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G137), .A2(new_n854), .B1(new_n800), .B2(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G159), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n798), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G143), .B2(new_n803), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n813), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n791), .A2(G132), .B1(G50), .B2(new_n809), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(new_n226), .C2(new_n769), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n781), .A2(new_n231), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n767), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n835), .A2(new_n821), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n767), .A2(new_n821), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n213), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n867), .A2(new_n763), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n848), .A2(new_n871), .ZN(G384));
  NOR2_X1   g0672(.A1(new_n694), .A2(new_n387), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n397), .B2(new_n399), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n375), .A2(new_n875), .A3(new_n388), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n375), .B2(new_n388), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n873), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n389), .B2(new_n400), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n744), .A2(new_n745), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n882), .A2(new_n883), .A3(new_n834), .ZN(new_n884));
  INV_X1    g0684(.A(new_n453), .ZN(new_n885));
  NOR2_X1   g0685(.A1(KEYINPUT104), .A2(KEYINPUT16), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n418), .B1(new_n812), .B2(new_n425), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n887), .A2(new_n231), .A3(new_n432), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n413), .ZN(new_n889));
  INV_X1    g0689(.A(new_n886), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n434), .A2(new_n414), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n293), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n437), .B1(new_n446), .B2(new_n445), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n689), .B1(new_n892), .B2(new_n437), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n885), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT105), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT105), .ZN(new_n898));
  INV_X1    g0698(.A(new_n894), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n453), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n898), .B(KEYINPUT37), .C1(new_n900), .C2(new_n893), .ZN(new_n901));
  INV_X1    g0701(.A(new_n689), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n438), .B1(new_n447), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n896), .A3(new_n453), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n455), .A2(new_n894), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n884), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n438), .A2(new_n902), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n450), .B2(new_n454), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n903), .A2(new_n453), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(new_n896), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n908), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n913), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n912), .A2(new_n913), .B1(new_n884), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(G330), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n403), .A2(new_n456), .A3(new_n458), .A4(new_n746), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n883), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n459), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n450), .A2(new_n902), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n389), .A2(KEYINPUT103), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n375), .A2(new_n875), .A3(new_n388), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n880), .B1(new_n929), .B2(new_n874), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n661), .B1(new_n504), .B2(new_n677), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n694), .B(new_n834), .C1(new_n931), .C2(new_n671), .ZN(new_n932));
  INV_X1    g0732(.A(new_n832), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n926), .B1(new_n934), .B2(new_n911), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n910), .A2(new_n918), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n929), .A2(new_n693), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n925), .B(new_n942), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n646), .B1(new_n459), .B2(new_n759), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n206), .B2(new_n684), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n571), .B1(new_n604), .B2(KEYINPUT35), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n947), .B(new_n241), .C1(KEYINPUT35), .C2(new_n604), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n242), .A2(new_n213), .A3(new_n410), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n201), .A2(new_n231), .ZN(new_n951));
  OAI211_X1 g0751(.A(G1), .B(new_n683), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n949), .A3(new_n952), .ZN(G367));
  INV_X1    g0753(.A(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n693), .A2(new_n611), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n631), .A3(new_n635), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n631), .A3(new_n958), .A4(new_n635), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n651), .A2(new_n694), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n954), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n954), .A3(new_n961), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n708), .A2(new_n703), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n677), .B1(new_n965), .B2(new_n709), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n970), .C1(new_n693), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n496), .A2(new_n498), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n659), .A3(new_n693), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n693), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n660), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT106), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n704), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n965), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n969), .A2(new_n970), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n971), .A2(new_n693), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n982), .B(new_n979), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n985), .ZN(new_n990));
  INV_X1    g0790(.A(new_n988), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n982), .B1(new_n972), .B2(new_n979), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n713), .B(KEYINPUT41), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n965), .A2(new_n710), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n965), .A2(KEYINPUT45), .A3(new_n710), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n965), .B2(new_n710), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n710), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1003), .A2(new_n963), .A3(KEYINPUT44), .A4(new_n964), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n981), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1000), .A2(new_n704), .A3(new_n1005), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n701), .A2(KEYINPUT109), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n708), .A2(new_n703), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n966), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n701), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1011), .B(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1007), .A2(new_n760), .A3(new_n1008), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n995), .B1(new_n1016), .B2(new_n760), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n989), .B(new_n993), .C1(new_n1017), .C2(new_n762), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n815), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n251), .B1(new_n210), .B2(new_n328), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n824), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n763), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT110), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n260), .B1(new_n777), .B2(new_n858), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n770), .A2(G68), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n783), .A2(new_n201), .B1(G58), .B2(new_n809), .ZN(new_n1026));
  INV_X1    g0826(.A(G143), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1026), .C1(new_n785), .C2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1024), .B(new_n1028), .C1(G77), .C2(new_n805), .ZN(new_n1029));
  INV_X1    g0829(.A(G137), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n791), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .C1(new_n283), .C2(new_n787), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n573), .A2(new_n798), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT111), .B(G311), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n854), .A2(new_n1035), .B1(G303), .B2(new_n803), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1034), .B(new_n1038), .C1(G294), .C2(new_n800), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n781), .A2(new_n215), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n814), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n789), .A2(new_n571), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT46), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1039), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n318), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n769), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1032), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT47), .Z(new_n1049));
  INV_X1    g0849(.A(new_n767), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1023), .B1(new_n978), .B2(new_n828), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1018), .A2(new_n1051), .ZN(G387));
  OR2_X1    g0852(.A1(new_n1015), .A2(new_n760), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1015), .A2(new_n760), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n713), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n703), .A2(new_n828), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n815), .B1(new_n248), .B2(new_n483), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n714), .B2(new_n819), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n715), .B1(G68), .B2(G77), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n324), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT50), .B1(new_n1060), .B2(G50), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1060), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n483), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1058), .A2(new_n1063), .B1(new_n228), .B2(new_n712), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n763), .B1(new_n1064), .B2(new_n1021), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n281), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n800), .A2(new_n1066), .B1(G50), .B2(new_n803), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n770), .A2(new_n327), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n283), .C2(new_n1031), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G77), .B2(new_n809), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n813), .B(new_n1040), .C1(new_n854), .C2(G159), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n231), .C2(new_n798), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT113), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n800), .A2(new_n1035), .B1(G303), .B2(new_n783), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1033), .B2(new_n787), .C1(new_n1075), .C2(new_n785), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT48), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n573), .B2(new_n769), .C1(new_n850), .C2(new_n789), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT49), .Z(new_n1079));
  OAI221_X1 g0879(.A(new_n813), .B1(new_n571), .B2(new_n781), .C1(new_n1031), .C2(new_n796), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1073), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1056), .B(new_n1065), .C1(new_n1081), .C2(new_n767), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n762), .B2(new_n1015), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1055), .A2(new_n1083), .ZN(G393));
  NAND3_X1  g0884(.A1(new_n1007), .A2(new_n762), .A3(new_n1008), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n963), .A2(new_n823), .A3(new_n964), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n785), .A2(new_n1033), .B1(new_n797), .B2(new_n787), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n769), .A2(new_n571), .B1(new_n573), .B2(new_n789), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n800), .B2(G303), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(new_n850), .C2(new_n798), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1031), .A2(new_n1075), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1091), .A2(new_n260), .A3(new_n782), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n800), .A2(new_n201), .B1(new_n324), .B2(new_n783), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n770), .A2(G77), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n231), .B2(new_n789), .C1(new_n221), .C2(new_n781), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n813), .B1(new_n1094), .B2(KEYINPUT114), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n785), .A2(new_n283), .B1(new_n858), .B2(new_n787), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G143), .B2(new_n791), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n767), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n824), .B1(new_n215), .B2(new_n210), .C1(new_n1019), .C2(new_n258), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1086), .A2(new_n763), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1085), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n720), .B1(new_n1108), .B2(new_n1054), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n1016), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  AND3_X1   g0911(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT38), .B1(new_n905), .B2(new_n906), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1112), .A2(new_n1113), .A3(new_n937), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n910), .B2(new_n918), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1114), .A2(new_n1115), .B1(new_n934), .B2(new_n940), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n940), .B1(new_n910), .B2(new_n918), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n833), .A2(new_n336), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n756), .A2(new_n694), .A3(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(new_n933), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n400), .A2(new_n879), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n927), .B2(new_n928), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1121), .B1(new_n1123), .B2(new_n880), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n878), .A2(new_n881), .A3(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1117), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1116), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n882), .A2(new_n834), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n841), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n930), .A2(new_n835), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n748), .B2(new_n749), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1116), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1131), .B1(new_n1137), .B2(new_n882), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n932), .A2(new_n933), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n746), .A2(new_n834), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n844), .A2(new_n1133), .B1(new_n1126), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1138), .A2(new_n1140), .B1(new_n1142), .B2(new_n1120), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n922), .B(new_n646), .C1(new_n459), .C2(new_n759), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1132), .B(new_n1136), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1126), .A2(new_n1141), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1134), .A2(new_n1147), .A3(new_n1120), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n834), .B1(new_n748), .B2(new_n749), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1149), .B2(new_n930), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1150), .B2(new_n1139), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1116), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1130), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1146), .B(new_n1151), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1145), .A2(new_n1154), .A3(new_n713), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT116), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1145), .A2(new_n1154), .A3(new_n1157), .A4(new_n713), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1139), .A2(new_n930), .B1(new_n693), .B2(new_n929), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n938), .A2(new_n939), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1119), .A2(new_n933), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1160), .A2(new_n1161), .B1(new_n1163), .B2(new_n1117), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1136), .B1(new_n1164), .B2(new_n1130), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n762), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n821), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n854), .A2(G128), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT54), .B(G143), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n783), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT53), .B1(new_n789), .B2(new_n283), .ZN(new_n1171));
  OR3_X1    g0971(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n283), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n769), .A2(new_n858), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n777), .A2(new_n1030), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n352), .B1(new_n805), .B2(new_n201), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n791), .A2(G125), .ZN(new_n1177));
  INV_X1    g0977(.A(G132), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1177), .C1(new_n1178), .C2(new_n787), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n800), .A2(new_n318), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n803), .A2(G116), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n783), .A2(G97), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1181), .A2(new_n1096), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1031), .A2(new_n850), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n785), .A2(new_n573), .ZN(new_n1186));
  OR3_X1    g0986(.A1(new_n865), .A2(new_n260), .A3(new_n790), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n767), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n281), .A2(new_n869), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1167), .A2(new_n763), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1159), .A2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(new_n869), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n201), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n299), .A2(new_n902), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n315), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n315), .A2(new_n1197), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OR3_X1    g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n763), .B1(new_n1204), .B2(new_n822), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1025), .B1(new_n777), .B2(new_n215), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n791), .A2(G283), .B1(G77), .B2(new_n809), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n805), .A2(G58), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1207), .A2(new_n267), .A3(new_n813), .A4(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT118), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1206), .B(new_n1210), .C1(new_n327), .C2(new_n783), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n228), .B2(new_n787), .C1(new_n571), .C2(new_n785), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT58), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G33), .A2(G41), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT117), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n218), .B(new_n1215), .C1(new_n814), .C2(G41), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n791), .B2(G124), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n858), .B2(new_n781), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n854), .A2(G125), .B1(new_n809), .B2(new_n1169), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n803), .A2(G128), .B1(G137), .B2(new_n783), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n283), .C2(new_n769), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G132), .B2(new_n800), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT59), .Z(new_n1223));
  OAI211_X1 g1023(.A(new_n1213), .B(new_n1216), .C1(new_n1218), .C2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1196), .B(new_n1205), .C1(new_n767), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1204), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n942), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n935), .A2(new_n941), .A3(new_n1204), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(G330), .A3(new_n920), .A4(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n935), .A2(new_n941), .A3(new_n1204), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1204), .B1(new_n935), .B2(new_n941), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n921), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1225), .B1(new_n1233), .B2(new_n762), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1154), .A2(new_n1146), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n713), .B1(new_n1235), .B2(KEYINPUT57), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1144), .B1(new_n1165), .B2(new_n1151), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1234), .B1(new_n1236), .B2(new_n1240), .ZN(G375));
  OAI21_X1  g1041(.A(new_n352), .B1(new_n789), .B2(new_n215), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n800), .A2(G116), .B1(G303), .B2(new_n791), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1068), .C1(new_n1046), .C2(new_n798), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(G77), .C2(new_n805), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n573), .B2(new_n787), .C1(new_n850), .C2(new_n785), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT119), .Z(new_n1247));
  OAI21_X1  g1047(.A(new_n814), .B1(new_n218), .B2(new_n769), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n800), .A2(new_n1169), .B1(G137), .B2(new_n803), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1178), .B2(new_n785), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT120), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n791), .A2(G128), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n783), .A2(G150), .B1(G159), .B2(new_n809), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1248), .B(new_n1256), .C1(G58), .C2(new_n805), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n767), .B1(new_n1247), .B2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1258), .B(new_n763), .C1(G68), .C2(new_n1195), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n821), .B2(new_n1126), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1151), .B2(new_n762), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1144), .B(new_n1148), .C1(new_n1150), .C2(new_n1139), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n994), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT121), .Z(G381));
  XOR2_X1   g1066(.A(G375), .B(KEYINPUT122), .Z(new_n1267));
  NAND2_X1  g1067(.A1(new_n1193), .A2(new_n1155), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1270), .A2(G384), .A3(G381), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1016), .A2(new_n760), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n762), .B1(new_n1273), .B2(new_n994), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n993), .A2(new_n989), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1051), .B(new_n1110), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1272), .A3(new_n1277), .ZN(G407));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  AND2_X1   g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1280), .A2(new_n1272), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1110), .B1(new_n1018), .B2(new_n1051), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1280), .A2(new_n1272), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1276), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT125), .B1(new_n1263), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1263), .A2(KEYINPUT125), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1289), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n713), .B(new_n1262), .C1(new_n1291), .C2(KEYINPUT60), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1261), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G384), .B(new_n1261), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n690), .A2(G213), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(G2897), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1298), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1235), .A2(new_n994), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1268), .B1(new_n1306), .B2(new_n1234), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT123), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1192), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(G375), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1235), .A2(KEYINPUT57), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1239), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n713), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(G378), .A2(KEYINPUT123), .A3(new_n1234), .A4(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1307), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1305), .B1(new_n1315), .B2(new_n1301), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1315), .A2(new_n1301), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1288), .B(new_n1316), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1307), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1317), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1300), .A3(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1287), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1287), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1316), .A2(new_n1288), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1330), .B1(new_n1318), .B2(KEYINPUT63), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1325), .A2(KEYINPUT126), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1318), .A2(KEYINPUT63), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1329), .A2(new_n1331), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1327), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1269), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1321), .A2(new_n1287), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1287), .B1(new_n1321), .B2(new_n1337), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT127), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1321), .A2(new_n1337), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1328), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT127), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1321), .A2(new_n1287), .A3(new_n1337), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1342), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1317), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1340), .A2(new_n1345), .A3(new_n1324), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


