

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595;

  XOR2_X1 U327 ( .A(n405), .B(KEYINPUT41), .Z(n576) );
  XOR2_X1 U328 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n357) );
  NOR2_X1 U329 ( .A1(n557), .A2(n531), .ZN(n431) );
  XNOR2_X1 U330 ( .A(n552), .B(KEYINPUT36), .ZN(n496) );
  XNOR2_X1 U331 ( .A(n414), .B(n413), .ZN(n557) );
  INV_X1 U332 ( .A(KEYINPUT79), .ZN(n372) );
  INV_X1 U333 ( .A(G204GAT), .ZN(n457) );
  XNOR2_X1 U334 ( .A(n568), .B(n372), .ZN(n552) );
  XNOR2_X1 U335 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U336 ( .A(n460), .B(n459), .ZN(G1353GAT) );
  XOR2_X1 U337 ( .A(G176GAT), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U338 ( .A(G43GAT), .B(G99GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U340 ( .A(G15GAT), .B(n297), .Z(n299) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U343 ( .A(G71GAT), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U344 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U346 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U347 ( .A(KEYINPUT0), .B(G127GAT), .Z(n305) );
  XNOR2_X1 U348 ( .A(KEYINPUT84), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U350 ( .A(G113GAT), .B(n306), .Z(n448) );
  XOR2_X1 U351 ( .A(KEYINPUT19), .B(G190GAT), .Z(n308) );
  XNOR2_X1 U352 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(n309), .ZN(n429) );
  XOR2_X1 U355 ( .A(n448), .B(n429), .Z(n310) );
  XOR2_X1 U356 ( .A(n311), .B(n310), .Z(n533) );
  INV_X1 U357 ( .A(n533), .ZN(n542) );
  XOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT21), .Z(n418) );
  XOR2_X1 U359 ( .A(G204GAT), .B(G148GAT), .Z(n383) );
  XOR2_X1 U360 ( .A(n418), .B(n383), .Z(n313) );
  XOR2_X1 U361 ( .A(G218GAT), .B(G162GAT), .Z(n353) );
  XOR2_X1 U362 ( .A(G155GAT), .B(G78GAT), .Z(n334) );
  XNOR2_X1 U363 ( .A(n353), .B(n334), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U365 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n315) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n432) );
  XOR2_X1 U368 ( .A(G22GAT), .B(n432), .Z(n317) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U372 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n321) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT24), .Z(n323) );
  XNOR2_X1 U376 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n474) );
  NOR2_X1 U380 ( .A1(n542), .A2(n474), .ZN(n328) );
  XOR2_X1 U381 ( .A(KEYINPUT26), .B(n328), .Z(n329) );
  XOR2_X1 U382 ( .A(KEYINPUT99), .B(n329), .Z(n476) );
  INV_X1 U383 ( .A(n476), .ZN(n555) );
  XOR2_X1 U384 ( .A(G1GAT), .B(KEYINPUT72), .Z(n331) );
  XNOR2_X1 U385 ( .A(G15GAT), .B(G22GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n392) );
  XNOR2_X1 U387 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n332), .B(KEYINPUT13), .ZN(n382) );
  XNOR2_X1 U389 ( .A(n392), .B(n382), .ZN(n347) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(G183GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n333), .B(G211GAT), .ZN(n426) );
  XOR2_X1 U392 ( .A(n426), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U393 ( .A(G127GAT), .B(n334), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n338) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U399 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n342) );
  XNOR2_X1 U400 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n343), .B(KEYINPUT81), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n347), .B(n346), .Z(n590) );
  INV_X1 U405 ( .A(n590), .ZN(n498) );
  XOR2_X1 U406 ( .A(G43GAT), .B(G29GAT), .Z(n349) );
  XNOR2_X1 U407 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(n350), .B(KEYINPUT71), .Z(n352) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n403) );
  XOR2_X1 U412 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n355) );
  XOR2_X1 U413 ( .A(G134GAT), .B(KEYINPUT78), .Z(n444) );
  XNOR2_X1 U414 ( .A(n353), .B(n444), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n361) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n359) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U421 ( .A1(n362), .A2(KEYINPUT66), .ZN(n366) );
  INV_X1 U422 ( .A(n362), .ZN(n364) );
  INV_X1 U423 ( .A(KEYINPUT66), .ZN(n363) );
  NAND2_X1 U424 ( .A1(n364), .A2(n363), .ZN(n365) );
  NAND2_X1 U425 ( .A1(n366), .A2(n365), .ZN(n370) );
  XOR2_X1 U426 ( .A(G92GAT), .B(G85GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G106GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U429 ( .A(G190GAT), .B(n381), .Z(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U431 ( .A(n403), .B(n371), .Z(n568) );
  NOR2_X1 U432 ( .A1(n498), .A2(n496), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT45), .ZN(n388) );
  XOR2_X1 U434 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n375) );
  XNOR2_X1 U435 ( .A(G120GAT), .B(G78GAT), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U437 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT75), .ZN(n377) );
  XOR2_X1 U439 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U440 ( .A1(G230GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n387) );
  XOR2_X1 U442 ( .A(n382), .B(n381), .Z(n385) );
  XOR2_X1 U443 ( .A(G176GAT), .B(G64GAT), .Z(n417) );
  XNOR2_X1 U444 ( .A(n383), .B(n417), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n468) );
  INV_X1 U447 ( .A(n468), .ZN(n405) );
  NAND2_X1 U448 ( .A1(n388), .A2(n405), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n389), .B(KEYINPUT115), .ZN(n404) );
  XOR2_X1 U450 ( .A(G169GAT), .B(G113GAT), .Z(n391) );
  NAND2_X1 U451 ( .A1(G229GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U453 ( .A(n393), .B(n392), .Z(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n395) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(G197GAT), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U457 ( .A(G8GAT), .B(KEYINPUT29), .Z(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U462 ( .A(n403), .B(n402), .Z(n517) );
  XOR2_X1 U463 ( .A(KEYINPUT73), .B(n517), .Z(n573) );
  NAND2_X1 U464 ( .A1(n404), .A2(n573), .ZN(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n410) );
  XOR2_X1 U466 ( .A(n590), .B(KEYINPUT113), .Z(n583) );
  NOR2_X1 U467 ( .A1(n517), .A2(n576), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n406), .B(KEYINPUT46), .ZN(n407) );
  NOR2_X1 U469 ( .A1(n583), .A2(n407), .ZN(n408) );
  NAND2_X1 U470 ( .A1(n408), .A2(n568), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U472 ( .A1(n412), .A2(n411), .ZN(n414) );
  XOR2_X1 U473 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n416) );
  XNOR2_X1 U475 ( .A(G36GAT), .B(G204GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n422) );
  XOR2_X1 U477 ( .A(G92GAT), .B(n417), .Z(n420) );
  XNOR2_X1 U478 ( .A(G218GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n425), .B(KEYINPUT95), .Z(n428) );
  XNOR2_X1 U484 ( .A(n426), .B(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n469) );
  BUF_X1 U487 ( .A(n469), .Z(n531) );
  XNOR2_X1 U488 ( .A(KEYINPUT54), .B(n431), .ZN(n453) );
  XOR2_X1 U489 ( .A(n432), .B(KEYINPUT89), .Z(n434) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n452) );
  XOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n436) );
  XNOR2_X1 U493 ( .A(G57GAT), .B(KEYINPUT90), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U495 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n438) );
  XNOR2_X1 U496 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U498 ( .A(n440), .B(n439), .Z(n450) );
  XOR2_X1 U499 ( .A(G85GAT), .B(G148GAT), .Z(n442) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(G162GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U502 ( .A(n444), .B(n443), .Z(n446) );
  XNOR2_X1 U503 ( .A(G29GAT), .B(G155GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n480) );
  INV_X1 U508 ( .A(n480), .ZN(n529) );
  NAND2_X1 U509 ( .A1(n453), .A2(n529), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT65), .ZN(n461) );
  NAND2_X1 U511 ( .A1(n555), .A2(n461), .ZN(n456) );
  INV_X1 U512 ( .A(KEYINPUT125), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n593) );
  INV_X1 U514 ( .A(n593), .ZN(n591) );
  NAND2_X1 U515 ( .A1(n591), .A2(n468), .ZN(n460) );
  XOR2_X1 U516 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n458) );
  NAND2_X1 U517 ( .A1(n474), .A2(n461), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT55), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n542), .ZN(n572) );
  NOR2_X1 U520 ( .A1(n552), .A2(n572), .ZN(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n465) );
  INV_X1 U522 ( .A(G190GAT), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  NOR2_X1 U525 ( .A1(n573), .A2(n468), .ZN(n503) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT27), .ZN(n477) );
  NOR2_X1 U527 ( .A1(n529), .A2(n477), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT97), .B(n470), .Z(n556) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT28), .ZN(n536) );
  NAND2_X1 U530 ( .A1(n556), .A2(n536), .ZN(n540) );
  XNOR2_X1 U531 ( .A(KEYINPUT98), .B(n540), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n542), .A2(n471), .ZN(n483) );
  NOR2_X1 U533 ( .A1(n531), .A2(n533), .ZN(n472) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(n472), .Z(n473) );
  NAND2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(KEYINPUT25), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n482) );
  NOR2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n497) );
  NAND2_X1 U541 ( .A1(n552), .A2(n590), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n484), .ZN(n485) );
  NOR2_X1 U543 ( .A1(n497), .A2(n485), .ZN(n518) );
  NAND2_X1 U544 ( .A1(n503), .A2(n518), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n529), .A2(n494), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(n486), .Z(n487) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U548 ( .A1(n531), .A2(n494), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n533), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n491) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT103), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n536), .A2(n494), .ZN(n495) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  NOR2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n499) );
  NAND2_X1 U559 ( .A1(n499), .A2(n498), .ZN(n502) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT104), .B(n500), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n527) );
  NAND2_X1 U563 ( .A1(n527), .A2(n503), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n504), .B(KEYINPUT38), .ZN(n505) );
  XNOR2_X1 U565 ( .A(KEYINPUT106), .B(n505), .ZN(n514) );
  NOR2_X1 U566 ( .A1(n529), .A2(n514), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n531), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n511) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n513) );
  NOR2_X1 U575 ( .A1(n533), .A2(n514), .ZN(n512) );
  XOR2_X1 U576 ( .A(n513), .B(n512), .Z(G1330GAT) );
  NOR2_X1 U577 ( .A1(n536), .A2(n514), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(n515), .Z(n516) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n516), .ZN(G1331GAT) );
  INV_X1 U580 ( .A(n517), .ZN(n585) );
  NOR2_X1 U581 ( .A1(n585), .A2(n576), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n528), .A2(n518), .ZN(n523) );
  NOR2_X1 U583 ( .A1(n529), .A2(n523), .ZN(n519) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(KEYINPUT42), .B(n520), .ZN(G1332GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n521), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n523), .ZN(n522) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n536), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(G78GAT), .B(n526), .Z(G1335GAT) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U595 ( .A1(n529), .A2(n535), .ZN(n530) );
  XOR2_X1 U596 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n535), .ZN(n532) );
  XOR2_X1 U598 ( .A(G92GAT), .B(n532), .Z(G1337GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U602 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(G106GAT), .B(n539), .Z(G1339GAT) );
  NOR2_X1 U605 ( .A1(n557), .A2(n540), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n573), .A2(n551), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(n543), .Z(n544) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  NOR2_X1 U610 ( .A1(n576), .A2(n551), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n549) );
  INV_X1 U614 ( .A(n551), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n547), .A2(n583), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  XOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT119), .Z(n561) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT118), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n570), .A2(n585), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1344GAT) );
  XNOR2_X1 U627 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n566) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  INV_X1 U629 ( .A(n576), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n562), .A2(n570), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n590), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U635 ( .A(n568), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1348GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n572), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n578) );
  XNOR2_X1 U643 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT56), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1349GAT) );
  INV_X1 U647 ( .A(n572), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n591), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G211GAT), .B(n592), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n496), .A2(n593), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

