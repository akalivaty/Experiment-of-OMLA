

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758;

  NOR2_X1 U378 ( .A1(n600), .A2(n528), .ZN(n529) );
  INV_X1 U379 ( .A(G953), .ZN(n399) );
  NOR2_X1 U380 ( .A1(n661), .A2(n675), .ZN(n603) );
  XOR2_X1 U381 ( .A(G125), .B(G146), .Z(n511) );
  NOR2_X1 U382 ( .A1(n567), .A2(n596), .ZN(n689) );
  XNOR2_X1 U383 ( .A(n529), .B(KEYINPUT0), .ZN(n571) );
  XNOR2_X1 U384 ( .A(n615), .B(KEYINPUT19), .ZN(n600) );
  AND2_X4 U385 ( .A1(n420), .A2(n358), .ZN(n725) );
  NOR2_X2 U386 ( .A1(n757), .A2(n758), .ZN(n384) );
  XNOR2_X2 U387 ( .A(n389), .B(KEYINPUT31), .ZN(n666) );
  NOR2_X2 U388 ( .A1(n454), .A2(n449), .ZN(n555) );
  NOR2_X2 U389 ( .A1(n557), .A2(n390), .ZN(n389) );
  INV_X1 U390 ( .A(n571), .ZN(n557) );
  XNOR2_X1 U391 ( .A(n511), .B(n470), .ZN(n744) );
  XNOR2_X1 U392 ( .A(G128), .B(KEYINPUT78), .ZN(n475) );
  NOR2_X1 U393 ( .A1(n709), .A2(G953), .ZN(n710) );
  XNOR2_X1 U394 ( .A(n382), .B(n381), .ZN(n638) );
  XNOR2_X1 U395 ( .A(n441), .B(n440), .ZN(n757) );
  NOR2_X1 U396 ( .A1(n557), .A2(n393), .ZN(n392) );
  XNOR2_X1 U397 ( .A(n426), .B(n507), .ZN(n596) );
  XNOR2_X1 U398 ( .A(n400), .B(n401), .ZN(n727) );
  XNOR2_X1 U399 ( .A(n402), .B(n404), .ZN(n400) );
  XNOR2_X1 U400 ( .A(n403), .B(n471), .ZN(n401) );
  XNOR2_X1 U401 ( .A(n477), .B(KEYINPUT3), .ZN(n516) );
  XNOR2_X1 U402 ( .A(n503), .B(KEYINPUT24), .ZN(n471) );
  XNOR2_X1 U403 ( .A(n475), .B(G143), .ZN(n513) );
  XNOR2_X1 U404 ( .A(G110), .B(G107), .ZN(n448) );
  XNOR2_X1 U405 ( .A(G119), .B(G113), .ZN(n477) );
  NOR2_X2 U406 ( .A1(n574), .A2(n647), .ZN(n576) );
  XNOR2_X2 U407 ( .A(n483), .B(n503), .ZN(n746) );
  INV_X1 U408 ( .A(G101), .ZN(n427) );
  XNOR2_X1 U409 ( .A(n384), .B(KEYINPUT46), .ZN(n383) );
  NOR2_X1 U410 ( .A1(n756), .A2(n655), .ZN(n584) );
  INV_X1 U411 ( .A(KEYINPUT103), .ZN(n436) );
  INV_X1 U412 ( .A(KEYINPUT4), .ZN(n428) );
  XOR2_X1 U413 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n501) );
  XNOR2_X1 U414 ( .A(KEYINPUT23), .B(KEYINPUT82), .ZN(n500) );
  XOR2_X1 U415 ( .A(G119), .B(G110), .Z(n505) );
  XNOR2_X1 U416 ( .A(n513), .B(n476), .ZN(n547) );
  INV_X1 U417 ( .A(G134), .ZN(n476) );
  XNOR2_X1 U418 ( .A(n499), .B(n498), .ZN(n545) );
  XNOR2_X1 U419 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n537) );
  XNOR2_X1 U421 ( .A(n534), .B(n433), .ZN(n536) );
  XNOR2_X1 U422 ( .A(n535), .B(n434), .ZN(n433) );
  INV_X1 U423 ( .A(G104), .ZN(n434) );
  XNOR2_X1 U424 ( .A(G122), .B(G113), .ZN(n530) );
  INV_X1 U425 ( .A(KEYINPUT10), .ZN(n470) );
  INV_X1 U426 ( .A(KEYINPUT48), .ZN(n381) );
  NAND2_X1 U427 ( .A1(n385), .A2(n383), .ZN(n382) );
  INV_X1 U428 ( .A(KEYINPUT44), .ZN(n419) );
  NAND2_X1 U429 ( .A1(G237), .A2(G234), .ZN(n523) );
  OR2_X1 U430 ( .A1(G902), .A2(G237), .ZN(n518) );
  AND2_X1 U431 ( .A1(n451), .A2(n604), .ZN(n450) );
  NAND2_X1 U432 ( .A1(n557), .A2(KEYINPUT34), .ZN(n451) );
  XNOR2_X1 U433 ( .A(n517), .B(n464), .ZN(n463) );
  XNOR2_X1 U434 ( .A(n513), .B(n465), .ZN(n464) );
  XNOR2_X1 U435 ( .A(n468), .B(KEYINPUT39), .ZN(n633) );
  NAND2_X1 U436 ( .A1(n395), .A2(n394), .ZN(n468) );
  NOR2_X1 U437 ( .A1(n357), .A2(n442), .ZN(n394) );
  INV_X1 U438 ( .A(n580), .ZN(n407) );
  NOR2_X1 U439 ( .A1(n618), .A2(n573), .ZN(n405) );
  XNOR2_X1 U440 ( .A(G478), .B(n553), .ZN(n566) );
  OR2_X1 U441 ( .A1(n727), .A2(G902), .ZN(n426) );
  INV_X1 U442 ( .A(KEYINPUT2), .ZN(n415) );
  NAND2_X1 U443 ( .A1(n399), .A2(G234), .ZN(n497) );
  XNOR2_X1 U444 ( .A(G140), .B(G143), .ZN(n535) );
  XNOR2_X1 U445 ( .A(n603), .B(n387), .ZN(n386) );
  INV_X1 U446 ( .A(KEYINPUT47), .ZN(n387) );
  AND2_X1 U447 ( .A1(n559), .A2(n455), .ZN(n453) );
  INV_X1 U448 ( .A(n557), .ZN(n559) );
  XOR2_X1 U449 ( .A(G137), .B(G131), .Z(n473) );
  XNOR2_X1 U450 ( .A(n414), .B(KEYINPUT74), .ZN(n413) );
  INV_X1 U451 ( .A(KEYINPUT5), .ZN(n414) );
  XNOR2_X1 U452 ( .A(n516), .B(n480), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n514), .B(KEYINPUT18), .ZN(n465) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT93), .Z(n510) );
  INV_X1 U455 ( .A(KEYINPUT68), .ZN(n447) );
  XNOR2_X1 U456 ( .A(n443), .B(n606), .ZN(n442) );
  AND2_X1 U457 ( .A1(n685), .A2(n594), .ZN(n595) );
  INV_X1 U458 ( .A(G469), .ZN(n487) );
  INV_X1 U459 ( .A(n690), .ZN(n461) );
  XNOR2_X1 U460 ( .A(n377), .B(n483), .ZN(n644) );
  XNOR2_X1 U461 ( .A(n378), .B(n485), .ZN(n377) );
  XNOR2_X1 U462 ( .A(n379), .B(n479), .ZN(n378) );
  XNOR2_X1 U463 ( .A(n478), .B(n413), .ZN(n479) );
  XNOR2_X1 U464 ( .A(n467), .B(n516), .ZN(n735) );
  XNOR2_X1 U465 ( .A(n546), .B(KEYINPUT16), .ZN(n467) );
  XOR2_X1 U466 ( .A(G140), .B(KEYINPUT67), .Z(n503) );
  XNOR2_X1 U467 ( .A(n506), .B(n502), .ZN(n404) );
  XNOR2_X1 U468 ( .A(G137), .B(G128), .ZN(n504) );
  XNOR2_X1 U469 ( .A(n539), .B(n435), .ZN(n720) );
  XNOR2_X1 U470 ( .A(n540), .B(n538), .ZN(n435) );
  INV_X1 U471 ( .A(KEYINPUT85), .ZN(n438) );
  XNOR2_X1 U472 ( .A(n509), .B(KEYINPUT69), .ZN(n429) );
  OR2_X1 U473 ( .A1(n614), .A2(n558), .ZN(n508) );
  INV_X1 U474 ( .A(KEYINPUT33), .ZN(n509) );
  XNOR2_X1 U475 ( .A(n667), .B(n432), .ZN(n632) );
  INV_X1 U476 ( .A(KEYINPUT110), .ZN(n432) );
  NAND2_X1 U477 ( .A1(n398), .A2(G953), .ZN(n591) );
  INV_X1 U478 ( .A(n590), .ZN(n398) );
  NAND2_X1 U479 ( .A1(n408), .A2(n406), .ZN(n376) );
  NOR2_X1 U480 ( .A1(n461), .A2(n375), .ZN(n370) );
  NAND2_X1 U481 ( .A1(n376), .A2(n372), .ZN(n371) );
  NOR2_X1 U482 ( .A1(n373), .A2(KEYINPUT88), .ZN(n372) );
  INV_X1 U483 ( .A(n461), .ZN(n373) );
  OR2_X1 U484 ( .A1(n732), .A2(G953), .ZN(n733) );
  AND2_X1 U485 ( .A1(n396), .A2(G953), .ZN(n525) );
  INV_X1 U486 ( .A(G898), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n550), .B(n431), .ZN(n723) );
  XNOR2_X1 U488 ( .A(n552), .B(n551), .ZN(n431) );
  INV_X1 U489 ( .A(KEYINPUT40), .ZN(n440) );
  XNOR2_X1 U490 ( .A(n616), .B(n430), .ZN(n617) );
  XNOR2_X1 U491 ( .A(KEYINPUT90), .B(KEYINPUT36), .ZN(n430) );
  NAND2_X1 U492 ( .A1(n407), .A2(n405), .ZN(n577) );
  XNOR2_X1 U493 ( .A(n392), .B(n391), .ZN(n650) );
  INV_X1 U494 ( .A(KEYINPUT102), .ZN(n391) );
  NAND2_X1 U495 ( .A1(n395), .A2(n688), .ZN(n393) );
  NOR2_X1 U496 ( .A1(n374), .A2(n368), .ZN(n647) );
  NOR2_X1 U497 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U498 ( .A1(n371), .A2(n369), .ZN(n368) );
  NOR2_X1 U499 ( .A1(n370), .A2(n596), .ZN(n369) );
  INV_X1 U500 ( .A(KEYINPUT56), .ZN(n457) );
  XNOR2_X1 U501 ( .A(n416), .B(KEYINPUT122), .ZN(n709) );
  AND2_X1 U502 ( .A1(n614), .A2(n462), .ZN(n355) );
  NOR2_X1 U503 ( .A1(n706), .A2(n361), .ZN(n356) );
  INV_X1 U504 ( .A(n624), .ZN(n594) );
  NAND2_X1 U505 ( .A1(n676), .A2(n594), .ZN(n357) );
  OR2_X1 U506 ( .A1(n732), .A2(n643), .ZN(n358) );
  NOR2_X1 U507 ( .A1(n607), .A2(n442), .ZN(n359) );
  OR2_X1 U508 ( .A1(n673), .A2(n732), .ZN(n360) );
  INV_X1 U509 ( .A(KEYINPUT34), .ZN(n455) );
  AND2_X1 U510 ( .A1(n708), .A2(n707), .ZN(n361) );
  INV_X1 U511 ( .A(KEYINPUT87), .ZN(n462) );
  XOR2_X1 U512 ( .A(G902), .B(KEYINPUT15), .Z(n635) );
  XOR2_X1 U513 ( .A(n711), .B(n712), .Z(n362) );
  XOR2_X1 U514 ( .A(n645), .B(KEYINPUT62), .Z(n363) );
  INV_X1 U515 ( .A(KEYINPUT88), .ZN(n375) );
  XOR2_X1 U516 ( .A(n720), .B(n719), .Z(n364) );
  XNOR2_X1 U517 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n365) );
  XNOR2_X1 U518 ( .A(KEYINPUT60), .B(KEYINPUT125), .ZN(n366) );
  AND2_X1 U519 ( .A1(n397), .A2(G953), .ZN(n729) );
  INV_X1 U520 ( .A(n729), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n512), .B(n367), .ZN(n515) );
  XNOR2_X2 U522 ( .A(n743), .B(n427), .ZN(n367) );
  XNOR2_X1 U523 ( .A(n367), .B(n380), .ZN(n485) );
  XNOR2_X1 U524 ( .A(n520), .B(n519), .ZN(n521) );
  NOR2_X1 U525 ( .A1(n684), .A2(n577), .ZN(n579) );
  NOR2_X2 U526 ( .A1(n732), .A2(n490), .ZN(n417) );
  INV_X1 U527 ( .A(G146), .ZN(n380) );
  NOR2_X1 U528 ( .A1(n388), .A2(n386), .ZN(n385) );
  NAND2_X1 U529 ( .A1(n619), .A2(n474), .ZN(n388) );
  NAND2_X1 U530 ( .A1(n650), .A2(n666), .ZN(n437) );
  INV_X1 U531 ( .A(n696), .ZN(n390) );
  INV_X1 U532 ( .A(n607), .ZN(n395) );
  NAND2_X1 U533 ( .A1(n359), .A2(n609), .ZN(n610) );
  NAND2_X1 U534 ( .A1(n399), .A2(G224), .ZN(n514) );
  AND2_X1 U535 ( .A1(n399), .A2(G227), .ZN(n472) );
  INV_X1 U536 ( .A(G952), .ZN(n397) );
  NAND2_X1 U537 ( .A1(n749), .A2(n399), .ZN(n754) );
  NAND2_X1 U538 ( .A1(n545), .A2(G221), .ZN(n402) );
  INV_X1 U539 ( .A(n744), .ZN(n403) );
  NAND2_X1 U540 ( .A1(n407), .A2(n355), .ZN(n406) );
  AND2_X1 U541 ( .A1(n410), .A2(n409), .ZN(n408) );
  OR2_X1 U542 ( .A1(n614), .A2(n462), .ZN(n409) );
  NAND2_X1 U543 ( .A1(n580), .A2(KEYINPUT87), .ZN(n410) );
  INV_X2 U544 ( .A(G122), .ZN(n411) );
  XNOR2_X2 U545 ( .A(n411), .B(G116), .ZN(n546) );
  NAND2_X1 U546 ( .A1(n412), .A2(n637), .ZN(n420) );
  NAND2_X1 U547 ( .A1(n417), .A2(n469), .ZN(n412) );
  NOR2_X1 U548 ( .A1(n688), .A2(n444), .ZN(n443) );
  XNOR2_X2 U549 ( .A(n481), .B(n482), .ZN(n688) );
  NAND2_X1 U550 ( .A1(n360), .A2(n415), .ZN(n446) );
  NAND2_X1 U551 ( .A1(n445), .A2(n356), .ZN(n416) );
  NAND2_X1 U552 ( .A1(n585), .A2(n418), .ZN(n586) );
  XNOR2_X1 U553 ( .A(n584), .B(n419), .ZN(n418) );
  XNOR2_X1 U554 ( .A(n460), .B(n362), .ZN(n459) );
  XNOR2_X1 U555 ( .A(n421), .B(n365), .ZN(G57) );
  NAND2_X1 U556 ( .A1(n425), .A2(n458), .ZN(n421) );
  XNOR2_X1 U557 ( .A(n422), .B(n366), .ZN(G60) );
  NAND2_X1 U558 ( .A1(n424), .A2(n458), .ZN(n422) );
  XNOR2_X1 U559 ( .A(n423), .B(n457), .ZN(G51) );
  NAND2_X1 U560 ( .A1(n459), .A2(n458), .ZN(n423) );
  XNOR2_X1 U561 ( .A(n721), .B(n364), .ZN(n424) );
  XNOR2_X1 U562 ( .A(n646), .B(n363), .ZN(n425) );
  XNOR2_X2 U563 ( .A(n572), .B(KEYINPUT22), .ZN(n580) );
  XNOR2_X1 U564 ( .A(n515), .B(n735), .ZN(n466) );
  XNOR2_X2 U565 ( .A(n428), .B(KEYINPUT65), .ZN(n743) );
  XNOR2_X2 U566 ( .A(n508), .B(n429), .ZN(n708) );
  XNOR2_X1 U567 ( .A(n673), .B(KEYINPUT75), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n466), .B(n463), .ZN(n711) );
  XNOR2_X1 U569 ( .A(n437), .B(n436), .ZN(n562) );
  XNOR2_X2 U570 ( .A(n439), .B(n438), .ZN(n673) );
  NAND2_X1 U571 ( .A1(n638), .A2(n634), .ZN(n439) );
  NAND2_X1 U572 ( .A1(n633), .A2(n625), .ZN(n441) );
  XNOR2_X2 U573 ( .A(n547), .B(n473), .ZN(n483) );
  INV_X1 U574 ( .A(n688), .ZN(n605) );
  INV_X1 U575 ( .A(n677), .ZN(n444) );
  NAND2_X1 U576 ( .A1(n446), .A2(n358), .ZN(n445) );
  XNOR2_X2 U577 ( .A(n736), .B(n447), .ZN(n517) );
  XNOR2_X2 U578 ( .A(n448), .B(G104), .ZN(n736) );
  NAND2_X1 U579 ( .A1(n452), .A2(n450), .ZN(n449) );
  NAND2_X1 U580 ( .A1(n708), .A2(n453), .ZN(n452) );
  NOR2_X1 U581 ( .A1(n708), .A2(n455), .ZN(n454) );
  XNOR2_X2 U582 ( .A(n517), .B(n472), .ZN(n484) );
  XNOR2_X2 U583 ( .A(n456), .B(KEYINPUT91), .ZN(n615) );
  NAND2_X1 U584 ( .A1(n608), .A2(n677), .ZN(n456) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n608) );
  NAND2_X1 U586 ( .A1(n725), .A2(G210), .ZN(n460) );
  XNOR2_X2 U587 ( .A(n589), .B(n588), .ZN(n732) );
  NOR2_X2 U588 ( .A1(G902), .A2(n713), .ZN(n488) );
  AND2_X1 U589 ( .A1(n598), .A2(n689), .ZN(n556) );
  XNOR2_X1 U590 ( .A(KEYINPUT81), .B(n660), .ZN(n474) );
  INV_X1 U591 ( .A(n669), .ZN(n619) );
  XNOR2_X1 U592 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U593 ( .A(n567), .ZN(n568) );
  INV_X1 U594 ( .A(KEYINPUT83), .ZN(n496) );
  AND2_X1 U595 ( .A1(n596), .A2(n595), .ZN(n612) );
  AND2_X1 U596 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U597 ( .A1(n622), .A2(n600), .ZN(n601) );
  XNOR2_X1 U598 ( .A(KEYINPUT70), .B(G472), .ZN(n482) );
  XNOR2_X1 U599 ( .A(G116), .B(KEYINPUT73), .ZN(n478) );
  NAND2_X1 U600 ( .A1(G210), .A2(n537), .ZN(n480) );
  NOR2_X1 U601 ( .A1(G902), .A2(n644), .ZN(n481) );
  XOR2_X1 U602 ( .A(n688), .B(KEYINPUT6), .Z(n614) );
  XOR2_X2 U603 ( .A(n485), .B(n484), .Z(n486) );
  XNOR2_X2 U604 ( .A(n486), .B(n746), .ZN(n713) );
  XNOR2_X2 U605 ( .A(n488), .B(n487), .ZN(n598) );
  XNOR2_X1 U606 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n489) );
  XNOR2_X2 U607 ( .A(n598), .B(n489), .ZN(n690) );
  INV_X1 U608 ( .A(n635), .ZN(n490) );
  NAND2_X1 U609 ( .A1(n490), .A2(G234), .ZN(n491) );
  XNOR2_X1 U610 ( .A(n491), .B(KEYINPUT20), .ZN(n493) );
  NAND2_X1 U611 ( .A1(G221), .A2(n493), .ZN(n492) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(n492), .Z(n685) );
  XOR2_X1 U613 ( .A(n685), .B(KEYINPUT100), .Z(n567) );
  XOR2_X1 U614 ( .A(KEYINPUT99), .B(KEYINPUT25), .Z(n495) );
  NAND2_X1 U615 ( .A1(n493), .A2(G217), .ZN(n494) );
  XNOR2_X1 U616 ( .A(n495), .B(n494), .ZN(n507) );
  XOR2_X1 U617 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n498) );
  XNOR2_X1 U618 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U619 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U620 ( .A1(n690), .A2(n689), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G214), .A2(n518), .ZN(n677) );
  NOR2_X1 U622 ( .A1(n635), .A2(n711), .ZN(n522) );
  NAND2_X1 U623 ( .A1(G210), .A2(n518), .ZN(n520) );
  XNOR2_X1 U624 ( .A(KEYINPUT95), .B(KEYINPUT79), .ZN(n519) );
  XOR2_X1 U625 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n524) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n526) );
  NAND2_X1 U627 ( .A1(n526), .A2(G952), .ZN(n705) );
  NOR2_X1 U628 ( .A1(G953), .A2(n705), .ZN(n593) );
  XOR2_X1 U629 ( .A(KEYINPUT96), .B(n525), .Z(n738) );
  NAND2_X1 U630 ( .A1(G902), .A2(n526), .ZN(n590) );
  NOR2_X1 U631 ( .A1(n738), .A2(n590), .ZN(n527) );
  NOR2_X1 U632 ( .A1(n593), .A2(n527), .ZN(n528) );
  XOR2_X1 U633 ( .A(KEYINPUT12), .B(KEYINPUT106), .Z(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(n530), .ZN(n540) );
  XOR2_X1 U635 ( .A(G131), .B(KEYINPUT11), .Z(n533) );
  XNOR2_X1 U636 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n532) );
  XNOR2_X1 U637 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U638 ( .A(n744), .B(n536), .Z(n539) );
  NAND2_X1 U639 ( .A1(n537), .A2(G214), .ZN(n538) );
  NOR2_X1 U640 ( .A1(n720), .A2(G902), .ZN(n544) );
  XOR2_X1 U641 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n542) );
  XNOR2_X1 U642 ( .A(KEYINPUT13), .B(G475), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n544), .B(n543), .ZN(n560) );
  INV_X1 U645 ( .A(n560), .ZN(n565) );
  NAND2_X1 U646 ( .A1(G217), .A2(n545), .ZN(n552) );
  XNOR2_X1 U647 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n551) );
  XOR2_X1 U648 ( .A(KEYINPUT109), .B(n546), .Z(n549) );
  XNOR2_X1 U649 ( .A(n547), .B(G107), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U651 ( .A1(G902), .A2(n723), .ZN(n553) );
  NOR2_X1 U652 ( .A1(n565), .A2(n566), .ZN(n604) );
  INV_X1 U653 ( .A(KEYINPUT35), .ZN(n554) );
  XNOR2_X1 U654 ( .A(n555), .B(n554), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n583), .A2(KEYINPUT44), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n556), .B(KEYINPUT101), .ZN(n607) );
  NOR2_X1 U657 ( .A1(n558), .A2(n688), .ZN(n696) );
  OR2_X1 U658 ( .A1(n566), .A2(n560), .ZN(n667) );
  NAND2_X1 U659 ( .A1(n566), .A2(n560), .ZN(n664) );
  INV_X1 U660 ( .A(n664), .ZN(n625) );
  NOR2_X1 U661 ( .A1(n632), .A2(n625), .ZN(n561) );
  XNOR2_X1 U662 ( .A(n561), .B(KEYINPUT111), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n562), .A2(n602), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n564), .A2(n563), .ZN(n574) );
  NAND2_X1 U665 ( .A1(n566), .A2(n565), .ZN(n678) );
  INV_X1 U666 ( .A(n678), .ZN(n569) );
  NAND2_X1 U667 ( .A1(n571), .A2(n570), .ZN(n572) );
  INV_X1 U668 ( .A(n614), .ZN(n573) );
  INV_X1 U669 ( .A(KEYINPUT89), .ZN(n575) );
  XNOR2_X1 U670 ( .A(n576), .B(n575), .ZN(n587) );
  INV_X1 U671 ( .A(n596), .ZN(n684) );
  XOR2_X1 U672 ( .A(KEYINPUT94), .B(n690), .Z(n618) );
  XNOR2_X1 U673 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n578) );
  XNOR2_X1 U674 ( .A(n579), .B(n578), .ZN(n756) );
  NOR2_X1 U675 ( .A1(n580), .A2(n690), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n688), .A2(n581), .ZN(n582) );
  NOR2_X1 U677 ( .A1(n684), .A2(n582), .ZN(n655) );
  BUF_X1 U678 ( .A(n583), .Z(n755) );
  NAND2_X1 U679 ( .A1(n584), .A2(n755), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n587), .A2(n586), .ZN(n589) );
  INV_X1 U681 ( .A(KEYINPUT45), .ZN(n588) );
  NOR2_X1 U682 ( .A1(G900), .A2(n591), .ZN(n592) );
  NOR2_X1 U683 ( .A1(n593), .A2(n592), .ZN(n624) );
  AND2_X1 U684 ( .A1(n605), .A2(n612), .ZN(n597) );
  XNOR2_X1 U685 ( .A(KEYINPUT28), .B(n597), .ZN(n599) );
  NAND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n622) );
  XNOR2_X1 U687 ( .A(n601), .B(KEYINPUT77), .ZN(n661) );
  INV_X1 U688 ( .A(n602), .ZN(n675) );
  INV_X1 U689 ( .A(n604), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n606) );
  INV_X1 U691 ( .A(n608), .ZN(n630) );
  NOR2_X1 U692 ( .A1(n624), .A2(n630), .ZN(n609) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n660) );
  NAND2_X1 U694 ( .A1(n625), .A2(n612), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n626), .A2(n615), .ZN(n616) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n669) );
  XNOR2_X1 U698 ( .A(KEYINPUT38), .B(KEYINPUT72), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(n630), .ZN(n676) );
  NAND2_X1 U700 ( .A1(n677), .A2(n676), .ZN(n674) );
  NOR2_X1 U701 ( .A1(n674), .A2(n678), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT41), .ZN(n699) );
  NOR2_X1 U703 ( .A1(n622), .A2(n699), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT42), .ZN(n758) );
  INV_X1 U705 ( .A(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n690), .A2(n627), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n628), .A2(n677), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT43), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n672) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n671) );
  AND2_X1 U711 ( .A1(n672), .A2(n671), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT84), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n672), .ZN(n641) );
  NAND2_X1 U715 ( .A1(KEYINPUT2), .A2(n671), .ZN(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT80), .B(n639), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U718 ( .A(KEYINPUT86), .B(n642), .Z(n643) );
  NAND2_X1 U719 ( .A1(n725), .A2(G472), .ZN(n646) );
  XOR2_X1 U720 ( .A(n644), .B(KEYINPUT113), .Z(n645) );
  XOR2_X1 U721 ( .A(n647), .B(G101), .Z(G3) );
  NOR2_X1 U722 ( .A1(n650), .A2(n664), .ZN(n648) );
  XOR2_X1 U723 ( .A(KEYINPUT114), .B(n648), .Z(n649) );
  XNOR2_X1 U724 ( .A(G104), .B(n649), .ZN(G6) );
  NOR2_X1 U725 ( .A1(n667), .A2(n650), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n652) );
  XNOR2_X1 U727 ( .A(G107), .B(KEYINPUT27), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(G9) );
  XOR2_X1 U730 ( .A(G110), .B(n655), .Z(G12) );
  NOR2_X1 U731 ( .A1(n661), .A2(n667), .ZN(n659) );
  XOR2_X1 U732 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n657) );
  XNOR2_X1 U733 ( .A(G128), .B(KEYINPUT116), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(G30) );
  XOR2_X1 U736 ( .A(G143), .B(n660), .Z(G45) );
  NOR2_X1 U737 ( .A1(n664), .A2(n661), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT118), .B(n662), .Z(n663) );
  XNOR2_X1 U739 ( .A(G146), .B(n663), .ZN(G48) );
  NOR2_X1 U740 ( .A1(n664), .A2(n666), .ZN(n665) );
  XOR2_X1 U741 ( .A(G113), .B(n665), .Z(G15) );
  NOR2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U743 ( .A(G116), .B(n668), .Z(G18) );
  XNOR2_X1 U744 ( .A(G125), .B(n669), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U746 ( .A(G134), .B(n671), .ZN(G36) );
  XNOR2_X1 U747 ( .A(G140), .B(n672), .ZN(G42) );
  NOR2_X1 U748 ( .A1(n675), .A2(n674), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n679) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n682), .B(KEYINPUT121), .ZN(n683) );
  NAND2_X1 U753 ( .A1(n683), .A2(n708), .ZN(n702) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT49), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT50), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT119), .B(n694), .Z(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT51), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(KEYINPUT120), .ZN(n700) );
  INV_X1 U764 ( .A(n699), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n700), .A2(n707), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U767 ( .A(KEYINPUT52), .B(n703), .Z(n704) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n710), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U770 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n712) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT123), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n725), .A2(G469), .ZN(n716) );
  XOR2_X1 U775 ( .A(n717), .B(n716), .Z(n718) );
  NOR2_X1 U776 ( .A1(n729), .A2(n718), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n725), .A2(G475), .ZN(n721) );
  XOR2_X1 U778 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n719) );
  NAND2_X1 U779 ( .A1(G478), .A2(n725), .ZN(n722) );
  XNOR2_X1 U780 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U781 ( .A1(n729), .A2(n724), .ZN(G63) );
  NAND2_X1 U782 ( .A1(G217), .A2(n725), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(G66) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U787 ( .A1(n731), .A2(G898), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(G101), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U792 ( .A(n741), .B(n740), .Z(n742) );
  XNOR2_X1 U793 ( .A(KEYINPUT126), .B(n742), .ZN(G69) );
  XNOR2_X1 U794 ( .A(KEYINPUT127), .B(n673), .ZN(n748) );
  XOR2_X1 U795 ( .A(n743), .B(n744), .Z(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n750) );
  INV_X1 U797 ( .A(n750), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U799 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U801 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U803 ( .A(G122), .B(n755), .Z(G24) );
  XOR2_X1 U804 ( .A(G119), .B(n756), .Z(G21) );
  XOR2_X1 U805 ( .A(n757), .B(G131), .Z(G33) );
  XOR2_X1 U806 ( .A(G137), .B(n758), .Z(G39) );
endmodule

