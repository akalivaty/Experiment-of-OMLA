//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT81), .B1(new_n193), .B2(G104), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n191), .A3(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n191), .A2(G107), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n193), .A2(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT5), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G116), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(G113), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G110), .B(G122), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n192), .A2(new_n194), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n197), .A2(new_n199), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT82), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n195), .A2(new_n222), .A3(new_n197), .A4(new_n199), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(G101), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n196), .A2(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  OR3_X1    g042(.A1(new_n214), .A2(KEYINPUT70), .A3(new_n206), .ZN(new_n229));
  INV_X1    g043(.A(new_n206), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n213), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n215), .A3(KEYINPUT70), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n217), .B(new_n218), .C1(new_n226), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT86), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n229), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n225), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n228), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT86), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n217), .A4(new_n218), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(G143), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G143), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n249), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n243), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(KEYINPUT65), .A3(new_n243), .A4(new_n258), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n253), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n256), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n268));
  INV_X1    g082(.A(new_n252), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n246), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT69), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT64), .B(G146), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n252), .B1(new_n274), .B2(G143), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n274), .B2(G143), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n273), .B(new_n275), .C1(new_n277), .C2(new_n265), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n267), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n264), .B1(new_n279), .B2(G125), .ZN(new_n280));
  INV_X1    g094(.A(G224), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n216), .B(new_n286), .C1(KEYINPUT88), .C2(new_n204), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n218), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT89), .B1(new_n205), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n212), .A2(new_n215), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n204), .B2(new_n286), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(new_n289), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n242), .A2(new_n285), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n280), .A2(new_n284), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT90), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT91), .B(new_n189), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n218), .B1(new_n239), .B2(new_n217), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT6), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n235), .B2(new_n241), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n302), .B2(new_n299), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n280), .B(new_n282), .Z(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n296), .B(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n294), .B1(new_n280), .B2(new_n284), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n241), .B2(new_n235), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT91), .B1(new_n311), .B2(new_n189), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n188), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n189), .B1(new_n295), .B2(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT91), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n187), .A3(new_n305), .A4(new_n298), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(KEYINPUT92), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n319), .B(new_n188), .C1(new_n306), .C2(new_n312), .ZN(new_n320));
  OAI21_X1  g134(.A(G214), .B1(G237), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(G122), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G122), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT14), .A3(G122), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G107), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT97), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT97), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(new_n332), .C1(KEYINPUT14), .C2(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n246), .A2(G128), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT95), .B1(new_n265), .B2(G143), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT95), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n246), .A3(G128), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n323), .A2(new_n325), .A3(new_n193), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT96), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n326), .A2(G107), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n345), .A2(new_n342), .B1(new_n339), .B2(new_n340), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT13), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT13), .B1(new_n336), .B2(new_n338), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(new_n348), .A3(new_n335), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT9), .B(G234), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(G217), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT98), .A3(new_n358), .ZN(new_n359));
  AOI211_X1 g173(.A(KEYINPUT98), .B(new_n357), .C1(new_n344), .C2(new_n350), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n361), .A3(new_n189), .ZN(new_n362));
  INV_X1    g176(.A(G478), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT15), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n362), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G113), .B(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(new_n191), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G125), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G140), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n274), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(KEYINPUT77), .A3(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n374), .B1(new_n378), .B2(new_n249), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n246), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT18), .A3(G131), .ZN(new_n385));
  INV_X1    g199(.A(new_n383), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n380), .B2(G214), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT93), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n379), .A2(new_n385), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n370), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  INV_X1    g214(.A(G131), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n388), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n384), .A2(G131), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n378), .B2(KEYINPUT19), .ZN(new_n405));
  OAI221_X1 g219(.A(new_n400), .B1(new_n402), .B2(new_n403), .C1(new_n405), .C2(new_n270), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n368), .B1(new_n395), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n249), .A3(new_n398), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n384), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n402), .A2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n410), .A2(KEYINPUT94), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n400), .A2(new_n414), .A3(new_n408), .A4(new_n409), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n413), .A2(new_n415), .B1(new_n394), .B2(new_n392), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n407), .B1(new_n416), .B2(new_n368), .ZN(new_n417));
  NOR2_X1   g231(.A1(G475), .A2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n415), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n368), .A3(new_n395), .ZN(new_n422));
  INV_X1    g236(.A(new_n407), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n418), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n421), .A2(new_n368), .A3(new_n395), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n368), .B1(new_n421), .B2(new_n395), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n189), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G475), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n366), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G952), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  INV_X1    g248(.A(G234), .ZN(new_n435));
  INV_X1    g249(.A(G237), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI211_X1 g252(.A(new_n189), .B(new_n354), .C1(G234), .C2(G237), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G898), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n432), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n318), .A2(new_n320), .A3(new_n321), .A4(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G469), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n256), .A2(new_n258), .A3(new_n266), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n265), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n256), .B2(new_n258), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n256), .A2(new_n258), .ZN(new_n450));
  INV_X1    g264(.A(new_n446), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n205), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n238), .A2(new_n263), .A3(new_n228), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n205), .A2(KEYINPUT10), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n456), .B(new_n457), .C1(new_n279), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G137), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT11), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n460), .A3(G134), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n462), .A2(new_n464), .B1(new_n340), .B2(G137), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(new_n401), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n354), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n272), .A2(new_n278), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n267), .B1(new_n200), .B2(new_n203), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n257), .B1(new_n274), .B2(G143), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT83), .B1(new_n477), .B2(new_n446), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n445), .A3(new_n452), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n475), .A2(new_n476), .B1(new_n479), .B2(new_n205), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n466), .B1(new_n480), .B2(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G128), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n273), .B1(new_n483), .B2(new_n275), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT69), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n454), .A3(KEYINPUT84), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n474), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT85), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n204), .A2(new_n445), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n278), .B2(new_n272), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n450), .A2(new_n451), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n267), .B1(new_n494), .B2(KEYINPUT83), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n204), .B1(new_n495), .B2(new_n452), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n491), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n466), .A3(new_n487), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n474), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n490), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n454), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n465), .B(G131), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(new_n474), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n473), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n459), .A2(new_n466), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n472), .B1(new_n468), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n444), .B(new_n189), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n444), .A2(new_n189), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n490), .A2(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n471), .B1(new_n512), .B2(new_n467), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n467), .A2(new_n471), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n509), .B(new_n511), .C1(new_n516), .C2(new_n444), .ZN(new_n517));
  INV_X1    g331(.A(G221), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n353), .B2(new_n189), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n443), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G217), .B1(new_n435), .B2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT73), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT24), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(G110), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G119), .B(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(G110), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT75), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n531), .A2(new_n538), .A3(new_n532), .A4(new_n535), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT76), .B1(new_n209), .B2(G128), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n540), .A2(KEYINPUT23), .B1(new_n209), .B2(G128), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(KEYINPUT23), .B2(new_n540), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n537), .A2(new_n539), .B1(G110), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n400), .A2(new_n408), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n531), .A2(new_n535), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n532), .A2(new_n546), .B1(new_n542), .B2(G110), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n399), .A2(G146), .B1(new_n274), .B2(new_n373), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n543), .A2(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT78), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n518), .A2(new_n435), .A3(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n552), .B2(new_n557), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n559), .A2(KEYINPUT25), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT25), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n525), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT79), .B(new_n525), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n550), .B2(new_n558), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n523), .A2(new_n189), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n263), .A2(new_n466), .ZN(new_n573));
  OR3_X1    g387(.A1(new_n460), .A2(KEYINPUT68), .A3(G134), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT68), .B1(new_n460), .B2(G134), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n461), .A3(new_n575), .ZN(new_n576));
  MUX2_X1   g390(.A(new_n576), .B(new_n465), .S(new_n401), .Z(new_n577));
  OAI211_X1 g391(.A(new_n573), .B(new_n236), .C1(new_n279), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n578), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT66), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n466), .B1(new_n263), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT66), .B(new_n253), .C1(new_n261), .C2(new_n262), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT67), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT65), .B1(new_n477), .B2(new_n243), .ZN(new_n586));
  INV_X1    g400(.A(new_n262), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n586), .A2(new_n587), .B1(new_n271), .B2(new_n245), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT66), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT67), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n263), .A2(new_n582), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n466), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n279), .A2(new_n577), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n585), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n581), .B1(new_n595), .B2(new_n237), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n580), .B1(new_n596), .B2(new_n579), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n380), .A2(G210), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT27), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT26), .B(G101), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n573), .B(KEYINPUT30), .C1(new_n279), .C2(new_n577), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n237), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT30), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n595), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n578), .A2(new_n601), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT31), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT71), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n607), .A2(KEYINPUT31), .A3(new_n608), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT71), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(KEYINPUT31), .C1(new_n607), .C2(new_n608), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n603), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT32), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n617), .A2(G472), .A3(G902), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n580), .B(new_n601), .C1(new_n596), .C2(new_n579), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n602), .B1(new_n607), .B2(new_n581), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT29), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT72), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n622), .B(new_n602), .C1(new_n578), .C2(new_n579), .ZN(new_n625));
  INV_X1    g439(.A(new_n573), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n237), .B1(new_n593), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n627), .A2(new_n578), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n624), .B(new_n625), .C1(new_n628), .C2(new_n579), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n579), .B1(new_n627), .B2(new_n578), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n580), .A2(KEYINPUT29), .A3(new_n601), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT72), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n614), .A2(new_n619), .B1(new_n634), .B2(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n572), .B1(new_n618), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n522), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n313), .A2(new_n317), .ZN(new_n639));
  INV_X1    g453(.A(new_n441), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  INV_X1    g455(.A(new_n358), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n357), .B1(new_n344), .B2(new_n350), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n641), .B1(new_n645), .B2(new_n360), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n358), .B1(new_n356), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT33), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n363), .A2(G902), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n651), .A2(new_n652), .B1(new_n363), .B2(new_n362), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n420), .A2(new_n426), .B1(new_n430), .B2(G475), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n639), .A2(new_n321), .A3(new_n640), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n657));
  INV_X1    g471(.A(new_n321), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n313), .B2(new_n317), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n640), .A4(new_n655), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n572), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n517), .A2(new_n663), .A3(new_n520), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n614), .A2(new_n189), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n616), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT101), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  INV_X1    g486(.A(new_n366), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n431), .A2(KEYINPUT102), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n430), .B2(G475), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n427), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n659), .A2(new_n640), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n668), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT35), .B(G107), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  AOI22_X1  g498(.A1(new_n665), .A2(G472), .B1(new_n615), .B2(new_n614), .ZN(new_n685));
  INV_X1    g499(.A(new_n551), .ZN(new_n686));
  INV_X1    g500(.A(new_n554), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n570), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n565), .A2(new_n566), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n565), .A2(new_n566), .A3(new_n695), .A4(new_n692), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n685), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n443), .A3(new_n521), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT37), .B(G110), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  NAND2_X1  g514(.A1(new_n614), .A2(new_n619), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n634), .A2(G472), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT32), .B1(new_n614), .B2(new_n615), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n694), .B(new_n696), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(G900), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n438), .B1(new_n439), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n677), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n659), .A2(new_n517), .A3(new_n708), .A4(new_n520), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n265), .ZN(G30));
  NAND2_X1  g525(.A1(new_n318), .A2(new_n320), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT38), .Z(new_n713));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n601), .B1(new_n607), .B2(new_n581), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n628), .B2(new_n602), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n614), .B2(new_n619), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n618), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n425), .B1(new_n424), .B2(new_n418), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT20), .B(new_n419), .C1(new_n422), .C2(new_n423), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n421), .A2(new_n395), .ZN(new_n723));
  INV_X1    g537(.A(new_n368), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n725), .B2(new_n422), .ZN(new_n726));
  INV_X1    g540(.A(G475), .ZN(new_n727));
  OAI22_X1  g541(.A1(new_n721), .A2(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n673), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n720), .A2(new_n658), .A3(new_n693), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n515), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n503), .B1(new_n502), .B2(new_n491), .ZN(new_n732));
  AOI211_X1 g546(.A(KEYINPUT85), .B(KEYINPUT12), .C1(new_n732), .C2(new_n487), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n499), .B1(new_n498), .B2(new_n474), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n505), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n468), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n731), .B1(new_n736), .B2(new_n471), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n510), .B1(new_n737), .B2(G469), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n519), .B1(new_n738), .B2(new_n509), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n707), .B(KEYINPUT39), .Z(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT40), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT40), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n713), .A2(new_n730), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G143), .ZN(G45));
  AOI21_X1  g559(.A(new_n642), .B1(KEYINPUT99), .B2(new_n643), .ZN(new_n746));
  INV_X1    g560(.A(new_n649), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n641), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT33), .B1(new_n359), .B2(new_n361), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n652), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n362), .A2(new_n363), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n707), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n728), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n658), .B(new_n754), .C1(new_n313), .C2(new_n317), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n694), .A2(new_n696), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n618), .A2(new_n635), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n739), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G146), .ZN(G48));
  AOI21_X1  g573(.A(new_n508), .B1(new_n735), .B2(new_n514), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n760), .B2(G902), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n509), .A3(new_n520), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n663), .C1(new_n704), .C2(new_n703), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n661), .B2(new_n657), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT41), .B(G113), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G15));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n679), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT105), .B(G116), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G18));
  NAND2_X1  g583(.A1(new_n694), .A2(new_n696), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n618), .B2(new_n635), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n762), .A2(new_n442), .A3(new_n659), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G119), .ZN(G21));
  NAND2_X1  g588(.A1(new_n639), .A2(new_n321), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n761), .A2(new_n509), .A3(new_n520), .A4(new_n640), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n776), .A3(new_n729), .ZN(new_n777));
  INV_X1    g591(.A(new_n580), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n602), .B1(new_n630), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n611), .A2(new_n609), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n615), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n666), .A2(new_n663), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G122), .ZN(G24));
  INV_X1    g598(.A(new_n754), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n762), .A2(new_n659), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n666), .A2(new_n693), .A3(new_n781), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT106), .B(G125), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G27));
  AOI21_X1  g604(.A(new_n658), .B1(new_n318), .B2(new_n320), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n636), .A2(new_n791), .A3(new_n739), .A4(new_n785), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  AND4_X1   g609(.A1(new_n636), .A2(new_n791), .A3(new_n739), .A4(new_n708), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n340), .ZN(G36));
  OR2_X1    g611(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(G469), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT107), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n511), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  INV_X1    g617(.A(new_n509), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n511), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n519), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n740), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n667), .A2(new_n693), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n654), .A2(new_n752), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT43), .Z(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n791), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n460), .ZN(G39));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n807), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n520), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n808), .B1(KEYINPUT109), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n791), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n757), .A3(new_n663), .A4(new_n754), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT110), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  NAND2_X1  g646(.A1(new_n433), .A2(new_n354), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT116), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n827), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n761), .A2(new_n509), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n519), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n782), .A2(new_n438), .A3(new_n813), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n828), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n762), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n713), .A2(new_n321), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT50), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n828), .A2(new_n437), .A3(new_n843), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(new_n813), .ZN(new_n847));
  INV_X1    g661(.A(new_n787), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n719), .A2(new_n572), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n654), .A3(new_n653), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n845), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n636), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n762), .A2(new_n659), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n434), .B1(new_n840), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n851), .B2(new_n655), .ZN(new_n859));
  INV_X1    g673(.A(new_n841), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n835), .B2(new_n837), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n853), .A2(KEYINPUT51), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n856), .B(new_n859), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n739), .A2(new_n685), .A3(new_n663), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n432), .B(KEYINPUT111), .C1(new_n654), .C2(new_n752), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT111), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n653), .B2(new_n654), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n441), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n321), .A3(new_n320), .A4(new_n318), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n865), .A2(new_n870), .B1(new_n763), .B2(new_n679), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n764), .A3(new_n698), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n637), .A2(new_n773), .A3(new_n783), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n673), .A2(new_n707), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n427), .C1(new_n674), .C2(new_n676), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n705), .A2(new_n875), .B1(new_n787), .B2(new_n754), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n828), .A2(new_n521), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n796), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n872), .A2(new_n794), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n565), .A2(new_n566), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT112), .A3(new_n692), .A4(new_n753), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n693), .B2(new_n707), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n658), .B(new_n729), .C1(new_n313), .C2(new_n317), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n739), .A3(new_n719), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n758), .A2(new_n887), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n705), .A2(new_n709), .B1(new_n786), .B2(new_n787), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT52), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n758), .A2(new_n887), .ZN(new_n892));
  INV_X1    g706(.A(new_n709), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n762), .A2(new_n659), .A3(new_n785), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n893), .A2(new_n771), .B1(new_n894), .B2(new_n848), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n879), .A2(new_n880), .A3(new_n890), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT113), .B1(new_n896), .B2(new_n890), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n895), .A3(new_n891), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT52), .B1(new_n888), .B2(new_n889), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n876), .A2(new_n877), .ZN(new_n904));
  INV_X1    g718(.A(new_n796), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n792), .A2(new_n793), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n792), .A2(new_n793), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n763), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n667), .A2(new_n770), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n662), .A2(new_n909), .B1(new_n522), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n318), .A2(new_n321), .A3(new_n320), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n432), .A2(KEYINPUT111), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n654), .A2(new_n752), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n640), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n909), .A2(new_n680), .B1(new_n668), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n772), .A2(new_n771), .B1(new_n777), .B2(new_n782), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n911), .A2(new_n918), .A3(new_n637), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n903), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT114), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n897), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n879), .B1(new_n898), .B2(new_n902), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT114), .B1(new_n926), .B2(KEYINPUT53), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(KEYINPUT53), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n879), .A2(new_n890), .A3(new_n896), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(KEYINPUT53), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n834), .B1(new_n864), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n713), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT49), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n836), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n836), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n520), .A2(new_n321), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n812), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n850), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n941), .ZN(G75));
  NOR2_X1   g756(.A1(new_n354), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  INV_X1    g759(.A(new_n897), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n921), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n923), .A3(new_n880), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n927), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G902), .ZN(new_n952));
  INV_X1    g766(.A(G210), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n303), .B(new_n304), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT55), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n944), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n956), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT117), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n954), .A2(KEYINPUT117), .A3(new_n956), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G51));
  XNOR2_X1  g776(.A(new_n510), .B(KEYINPUT57), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n925), .B1(new_n924), .B2(new_n927), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n506), .B2(new_n508), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n952), .A2(new_n801), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n943), .B1(new_n967), .B2(new_n968), .ZN(G54));
  NAND4_X1  g783(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n970), .A2(new_n417), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n417), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n943), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n928), .B2(new_n932), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n651), .B(KEYINPUT118), .Z(new_n977));
  OAI21_X1  g791(.A(new_n944), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n975), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n964), .B2(new_n965), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT119), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(KEYINPUT119), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT60), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n568), .B1(new_n951), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT121), .B1(new_n988), .B2(new_n943), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT121), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n924), .B2(new_n927), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n990), .B(new_n944), .C1(new_n991), .C2(new_n568), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n690), .B2(new_n691), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n988), .A2(new_n943), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(KEYINPUT61), .A3(new_n993), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(G66));
  OAI21_X1  g813(.A(G953), .B1(new_n440), .B2(new_n281), .ZN(new_n1000));
  INV_X1    g814(.A(new_n920), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(new_n303), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(G898), .B2(new_n354), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1002), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(new_n595), .A2(new_n606), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n604), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(new_n405), .Z(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT122), .Z(new_n1009));
  AND2_X1   g823(.A1(new_n895), .A2(new_n758), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n744), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT62), .Z(new_n1012));
  NAND2_X1  g826(.A1(new_n831), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT123), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n741), .B1(new_n868), .B2(new_n866), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1015), .A2(new_n636), .A3(new_n791), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1014), .B(new_n1016), .C1(new_n809), .C2(new_n818), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n809), .B2(new_n818), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT123), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1013), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1009), .B1(new_n1020), .B2(G953), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n354), .B1(G227), .B2(G900), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT124), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1010), .A2(new_n794), .A3(new_n905), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n819), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n808), .A2(new_n636), .A3(new_n740), .A4(new_n886), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1027), .A2(new_n354), .A3(new_n831), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1008), .B1(G900), .B2(G953), .ZN(new_n1030));
  AOI22_X1  g844(.A1(new_n1029), .A2(new_n1030), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1021), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1025), .B1(new_n1021), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1032), .A2(new_n1033), .ZN(G72));
  XNOR2_X1  g848(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n714), .A2(new_n189), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1035), .B(new_n1036), .Z(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  OR3_X1    g852(.A1(new_n607), .A2(new_n581), .A3(new_n601), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n931), .A2(new_n715), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1037), .B1(new_n1020), .B2(new_n1001), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1040), .B1(new_n1041), .B2(new_n715), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1039), .B(KEYINPUT126), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1027), .A2(new_n831), .A3(new_n1001), .A4(new_n1028), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n1045), .B2(new_n1038), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT127), .ZN(new_n1047));
  OR3_X1    g861(.A1(new_n1046), .A2(new_n1047), .A3(new_n943), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1047), .B1(new_n1046), .B2(new_n943), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(G57));
endmodule


