//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT68), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT69), .Z(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT70), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n471), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n486));
  INV_X1    g061(.A(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n487), .A2(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n490), .A2(new_n493), .B1(G102), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n488), .B2(new_n489), .ZN(new_n497));
  AND2_X1   g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n492), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(KEYINPUT71), .C1(new_n463), .C2(new_n462), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n491), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT73), .B1(new_n509), .B2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT73), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(KEYINPUT72), .A3(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT75), .B(G88), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n524), .B(new_n525), .C1(new_n517), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  INV_X1    g104(.A(new_n515), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n520), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT77), .B(G51), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n532), .A2(G543), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n536), .A2(KEYINPUT78), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT78), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT7), .Z(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT79), .B(G89), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n522), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  OAI21_X1  g121(.A(G543), .B1(new_n520), .B2(new_n533), .ZN(new_n547));
  AOI211_X1 g122(.A(KEYINPUT76), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n517), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT80), .B(G90), .Z(new_n553));
  NAND2_X1  g128(.A1(new_n522), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  NOR3_X1   g132(.A1(new_n547), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n513), .A2(new_n520), .A3(G81), .ZN(new_n559));
  AND2_X1   g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n513), .B2(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n561), .B2(new_n517), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT81), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n508), .B(new_n572), .C1(new_n510), .C2(new_n512), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT83), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n579), .B(G651), .C1(new_n574), .C2(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n582));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT9), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n549), .A2(new_n585), .A3(G53), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n584), .A2(new_n586), .B1(G91), .B2(new_n522), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n587), .ZN(G299));
  OAI21_X1  g163(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(G87), .ZN(new_n590));
  INV_X1    g165(.A(G49), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n590), .B2(new_n521), .C1(new_n582), .C2(new_n591), .ZN(G288));
  AOI22_X1  g167(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n517), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n520), .A2(G48), .A3(G543), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n521), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n513), .A2(G60), .ZN(new_n600));
  INV_X1    g175(.A(G72), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n507), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n522), .B2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n549), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n521), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n513), .A2(new_n520), .A3(new_n609), .A4(G92), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(KEYINPUT10), .B1(new_n608), .B2(new_n610), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n571), .B2(new_n573), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT85), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n549), .A2(G54), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT86), .B1(new_n620), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n606), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n606), .B1(new_n625), .B2(G868), .ZN(G321));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G168), .B2(new_n628), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(G168), .B2(new_n628), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n474), .A2(new_n494), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n476), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n479), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n642), .A2(new_n643), .A3(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT14), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(new_n666), .A3(G14), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  XOR2_X1   g247(.A(new_n670), .B(KEYINPUT88), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT17), .ZN(new_n674));
  INV_X1    g249(.A(new_n668), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n670), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n669), .B1(new_n678), .B2(KEYINPUT87), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(KEYINPUT87), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n674), .B2(new_n669), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(new_n649), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n677), .A2(new_n682), .A3(G2096), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n684), .A2(new_n641), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n641), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n692), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n690), .B1(new_n697), .B2(KEYINPUT89), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(KEYINPUT89), .B2(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT90), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  INV_X1    g281(.A(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n704), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n708), .B1(new_n705), .B2(new_n709), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G6), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n598), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT32), .B(G1981), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n713), .A2(G23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G288), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT91), .B(G16), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n724), .B(new_n725), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT34), .B1(new_n720), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n718), .B2(new_n719), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n476), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n479), .A2(G119), .ZN(new_n742));
  OR2_X1    g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(new_n739), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  XOR2_X1   g323(.A(new_n747), .B(new_n748), .Z(new_n749));
  NOR2_X1   g324(.A1(new_n727), .A2(G24), .ZN(new_n750));
  INV_X1    g325(.A(G290), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n727), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G1986), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(G1986), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n735), .A2(new_n738), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(KEYINPUT36), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n735), .A2(new_n738), .A3(new_n758), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n713), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n713), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G1966), .ZN(new_n764));
  NOR2_X1   g339(.A1(G5), .A2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G301), .B2(new_n713), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n648), .A2(new_n739), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n739), .B1(new_n772), .B2(G28), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n774), .B1(new_n772), .B2(G28), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n763), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n739), .A2(G32), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  INV_X1    g358(.A(G129), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n478), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n494), .A2(G105), .ZN(new_n786));
  INV_X1    g361(.A(G141), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n475), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(new_n739), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n739), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n799));
  OAI221_X1 g374(.A(G2104), .B1(G116), .B2(new_n471), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G140), .ZN(new_n801));
  INV_X1    g376(.A(G128), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n800), .B1(new_n475), .B2(new_n801), .C1(new_n802), .C2(new_n478), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n796), .B1(new_n804), .B2(new_n739), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT95), .B(G2067), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT24), .ZN(new_n809));
  INV_X1    g384(.A(G34), .ZN(new_n810));
  AOI21_X1  g385(.A(G29), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G160), .B2(new_n739), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n807), .B(new_n808), .C1(G2084), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n739), .A2(G27), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n739), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2078), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n794), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n726), .A2(G20), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G299), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1956), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n727), .A2(G19), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n563), .B2(new_n727), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1341), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n739), .A2(G35), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G162), .B2(new_n739), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT29), .B(G2090), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n790), .B2(new_n792), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n739), .A2(G33), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT25), .ZN(new_n836));
  NAND2_X1  g411(.A1(G115), .A2(G2104), .ZN(new_n837));
  INV_X1    g412(.A(G127), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n464), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(G2105), .ZN(new_n840));
  AOI211_X1 g415(.A(new_n836), .B(new_n840), .C1(G139), .C2(new_n476), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n834), .B1(new_n841), .B2(new_n739), .ZN(new_n842));
  INV_X1    g417(.A(G2072), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n767), .A2(new_n768), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n829), .A2(new_n831), .B1(G2084), .B2(new_n813), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n833), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR4_X1   g422(.A1(new_n818), .A2(new_n824), .A3(new_n827), .A4(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n763), .A2(new_n849), .A3(new_n764), .A4(new_n778), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n713), .A2(G4), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n625), .B2(new_n713), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT93), .B(G1348), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AND4_X1   g429(.A1(new_n780), .A2(new_n848), .A3(new_n850), .A4(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n760), .A2(new_n855), .ZN(G311));
  AND3_X1   g431(.A1(new_n760), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT101), .B1(new_n760), .B2(new_n855), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(G150));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n558), .B2(new_n562), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT102), .B(G55), .Z(new_n862));
  NAND4_X1  g437(.A1(new_n532), .A2(G543), .A3(new_n534), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n513), .A2(new_n520), .A3(G93), .ZN(new_n864));
  AND2_X1   g439(.A1(G80), .A2(G543), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n513), .B2(G67), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n517), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n532), .A2(G43), .A3(G543), .A4(new_n534), .ZN(new_n868));
  INV_X1    g443(.A(G56), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n505), .B1(new_n507), .B2(KEYINPUT74), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(KEYINPUT5), .A3(new_n511), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(new_n508), .ZN(new_n872));
  OAI21_X1  g447(.A(G651), .B1(new_n872), .B2(new_n560), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n868), .A2(new_n873), .A3(KEYINPUT103), .A4(new_n559), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n861), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n862), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n547), .A2(new_n548), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n864), .B1(new_n866), .B2(new_n517), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n563), .A2(new_n879), .A3(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT38), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n624), .A2(new_n632), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n882), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT104), .ZN(new_n888));
  AOI21_X1  g463(.A(G860), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n867), .A2(G860), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT37), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  XNOR2_X1  g468(.A(new_n803), .B(new_n503), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n841), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n789), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n789), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  OR2_X1    g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n899), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n900));
  INV_X1    g475(.A(G142), .ZN(new_n901));
  INV_X1    g476(.A(G130), .ZN(new_n902));
  OAI221_X1 g477(.A(new_n900), .B1(new_n475), .B2(new_n901), .C1(new_n902), .C2(new_n478), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n639), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(new_n746), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n746), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(new_n897), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n898), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(KEYINPUT105), .A3(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n648), .B(G160), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n483), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT107), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n909), .A2(new_n911), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n913), .A2(new_n897), .A3(new_n896), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(new_n916), .ZN(new_n924));
  AOI211_X1 g499(.A(KEYINPUT106), .B(new_n924), .C1(new_n920), .C2(new_n921), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n918), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g502(.A1(new_n634), .A2(new_n881), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n625), .A2(new_n632), .A3(new_n880), .A4(new_n875), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n522), .A2(G91), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n585), .B1(new_n549), .B2(G53), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT9), .A4(new_n583), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n578), .B2(new_n580), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n624), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT86), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n572), .B1(new_n871), .B2(new_n508), .ZN(new_n938));
  INV_X1    g513(.A(new_n573), .ZN(new_n939));
  OAI21_X1  g514(.A(G66), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n517), .B1(new_n940), .B2(new_n618), .ZN(new_n941));
  INV_X1    g516(.A(G54), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n582), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n937), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n621), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(G299), .A2(new_n946), .A3(new_n614), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n936), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n936), .A2(new_n947), .A3(KEYINPUT108), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n930), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT41), .B1(new_n936), .B2(new_n947), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n929), .B(new_n928), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  INV_X1    g532(.A(G288), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n751), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G290), .A2(G288), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(G305), .B(G303), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n957), .A3(new_n960), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n951), .A2(new_n969), .A3(new_n954), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n956), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n956), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(G868), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(G868), .B2(new_n879), .ZN(G295));
  OAI21_X1  g549(.A(new_n973), .B1(G868), .B2(new_n879), .ZN(G331));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT110), .A4(new_n554), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n544), .C1(new_n538), .C2(new_n539), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g555(.A1(G301), .A2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n875), .A2(new_n981), .A3(new_n880), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n875), .B2(new_n880), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n881), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n979), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n875), .A2(new_n981), .A3(new_n880), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n952), .B2(new_n953), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n936), .A2(new_n947), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n984), .A3(new_n989), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n968), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G37), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n949), .A2(new_n950), .A3(new_n989), .A4(new_n984), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n968), .B1(new_n997), .B2(new_n991), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n977), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n947), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n990), .A2(new_n1000), .A3(new_n948), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT41), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n992), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n936), .A2(new_n947), .A3(KEYINPUT41), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1003), .A2(new_n1004), .B1(new_n989), .B2(new_n984), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n967), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1006), .A2(KEYINPUT111), .A3(new_n995), .A4(new_n994), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n976), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n996), .ZN(new_n1009));
  INV_X1    g584(.A(new_n993), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n967), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT43), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n976), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n996), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(G397));
  NAND2_X1  g593(.A1(G286), .A2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT124), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1025), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1029), .B2(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n503), .A2(new_n1025), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1028), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT118), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1031), .B2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n503), .A2(new_n1041), .A3(new_n1025), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT119), .B(G2084), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1023), .B1(new_n1039), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1022), .B1(new_n1047), .B2(new_n1021), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1030), .A2(new_n1038), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n1023), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1038), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT118), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1019), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT124), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1048), .B1(new_n1058), .B2(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT62), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1047), .A2(KEYINPUT123), .B1(new_n1056), .B2(KEYINPUT124), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1021), .B1(new_n1064), .B2(new_n1051), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1063), .B(new_n1060), .C1(new_n1065), .C2(new_n1048), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT55), .B1(G166), .B2(new_n1023), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n1068));
  NAND3_X1  g643(.A1(G303), .A2(new_n1068), .A3(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1035), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n730), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1043), .A2(G2090), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1023), .B(new_n1070), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1070), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n503), .A2(KEYINPUT117), .A3(new_n1041), .A4(new_n1025), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1042), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1040), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(G2090), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1031), .A2(new_n1028), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n1023), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(G288), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n1087), .C1(new_n1088), .C2(G288), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n598), .A2(new_n707), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n1094));
  OAI21_X1  g669(.A(G1981), .B1(new_n594), .B2(new_n597), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n1097));
  NAND3_X1  g672(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1087), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1097), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1090), .B(new_n1092), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1077), .A2(new_n1085), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G2078), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT53), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1044), .A2(G1961), .B1(new_n1036), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1073), .B1(new_n1072), .B2(new_n1035), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G301), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1103), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1062), .A2(new_n1066), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n1111), .B2(G301), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1111), .B2(G301), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n1119), .B2(new_n1104), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(G171), .C1(new_n1120), .C2(new_n1106), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1120), .A2(G171), .A3(new_n1106), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1116), .B1(new_n1112), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1122), .A2(new_n1124), .A3(new_n1103), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1060), .B1(new_n1065), .B2(new_n1048), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G299), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1082), .A2(new_n823), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n581), .A2(new_n587), .A3(new_n1127), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1029), .A2(KEYINPUT121), .A3(new_n1130), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1129), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G2067), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1043), .A2(new_n853), .B1(new_n1137), .B2(new_n1086), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n624), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1138), .B(new_n624), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1145), .A2(KEYINPUT60), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT58), .B(G1341), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1036), .A2(G1996), .B1(new_n1086), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n563), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1152));
  NOR2_X1   g727(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n563), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1144), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1125), .A2(new_n1126), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1102), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1050), .A2(new_n1023), .A3(G286), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1078), .B1(new_n1164), .B2(G8), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT63), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n958), .A2(new_n1088), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1093), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1085), .A2(KEYINPUT63), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1077), .B1(new_n1173), .B2(new_n1162), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1102), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1114), .A2(new_n1160), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1033), .A2(new_n1028), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(KEYINPUT112), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(KEYINPUT112), .B2(new_n1180), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1178), .A2(G1986), .A3(G290), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT113), .Z(new_n1185));
  XNOR2_X1  g760(.A(new_n789), .B(G1996), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n803), .B(new_n1137), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n745), .B(new_n748), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1179), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1177), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1179), .B1(new_n1187), .B2(new_n789), .ZN(new_n1194));
  INV_X1    g769(.A(G1996), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1178), .A2(KEYINPUT46), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT46), .B1(new_n1178), .B2(new_n1195), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  INV_X1    g774(.A(KEYINPUT48), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1191), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1200), .B2(new_n1182), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n746), .A2(new_n748), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1188), .A2(new_n1203), .B1(G2067), .B2(new_n803), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1178), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1199), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1193), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g782(.A1(new_n710), .A2(new_n711), .A3(G401), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n686), .A2(G319), .A3(new_n687), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g787(.A1(new_n686), .A2(KEYINPUT126), .A3(G319), .A4(new_n687), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AND3_X1   g789(.A1(new_n1209), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1210), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n926), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1218), .A2(new_n1219), .ZN(G308));
  OAI221_X1 g794(.A(new_n926), .B1(new_n1015), .B2(new_n1016), .C1(new_n1217), .C2(new_n1216), .ZN(G225));
endmodule


