//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n210), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n210), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n206), .C2(new_n218), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(new_n233));
  NAND4_X1  g0033(.A1(new_n233), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n219), .A2(KEYINPUT0), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n220), .A2(new_n231), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT69), .B(G50), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT70), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n253), .B(new_n257), .ZN(G351));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n262), .B(new_n263), .C1(G1), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT85), .B1(new_n263), .B2(G97), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n263), .A2(KEYINPUT85), .A3(G97), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n266), .A2(G97), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT83), .ZN(new_n270));
  AND2_X1   g0070(.A1(G97), .A2(G107), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G97), .A2(G107), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT82), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(KEYINPUT6), .ZN(new_n274));
  MUX2_X1   g0074(.A(new_n273), .B(G97), .S(KEYINPUT6), .Z(new_n275));
  NAND2_X1  g0075(.A1(G97), .A2(G107), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n207), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n270), .B(new_n274), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n273), .A2(KEYINPUT6), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT6), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G97), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n207), .B(new_n276), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n270), .B1(new_n283), .B2(new_n274), .ZN(new_n284));
  OAI21_X1  g0084(.A(G20), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT7), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(KEYINPUT79), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT79), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n295), .B2(new_n264), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n286), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G107), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G77), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n285), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT84), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n303), .A2(new_n304), .A3(new_n261), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n303), .B2(new_n261), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n269), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n260), .B1(G33), .B2(G41), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G283), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n287), .A2(G1698), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n311), .C1(new_n210), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n228), .A2(G1698), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT4), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n308), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n211), .A2(G45), .ZN(new_n321));
  OR2_X1    g0121(.A1(KEYINPUT5), .A2(G41), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT5), .A2(G41), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n308), .ZN(new_n325));
  INV_X1    g0125(.A(G274), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n308), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n325), .A2(G257), .B1(new_n327), .B2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G169), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n307), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT10), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n308), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G41), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G1), .A3(G13), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n335), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(G226), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n287), .A2(G222), .A3(new_n309), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n227), .B2(new_n287), .C1(new_n312), .C2(new_n343), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n336), .B(new_n341), .C1(new_n344), .C2(new_n308), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n334), .B1(new_n347), .B2(KEYINPUT74), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n349), .A2(new_n250), .A3(KEYINPUT8), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(KEYINPUT71), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n212), .A3(G33), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n301), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n262), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n263), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n202), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n262), .B1(G1), .B2(new_n212), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n202), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n345), .A2(G190), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n347), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n348), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n348), .A2(new_n364), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n345), .A2(G169), .B1(new_n355), .B2(new_n359), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n345), .A2(new_n331), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n339), .A2(new_n228), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n371), .A2(new_n336), .A3(KEYINPUT72), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n312), .A2(new_n223), .B1(new_n206), .B2(new_n287), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n314), .A2(new_n290), .ZN(new_n374));
  INV_X1    g0174(.A(G232), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n374), .A2(new_n375), .A3(G1698), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n308), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT72), .B1(new_n371), .B2(new_n336), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n301), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n351), .A2(new_n382), .B1(new_n212), .B2(new_n227), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n212), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n261), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n356), .A2(new_n227), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n227), .C2(new_n358), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n381), .B(new_n389), .C1(G179), .C2(new_n379), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n389), .B(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n379), .A2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n379), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n367), .A2(new_n370), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n352), .A2(new_n356), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n358), .B2(new_n352), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n250), .A2(new_n222), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n201), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n301), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n299), .B2(G68), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n261), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n292), .A2(new_n294), .A3(G33), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n314), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n222), .B1(new_n409), .B2(new_n286), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT7), .B1(new_n317), .B2(G20), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n407), .B(new_n402), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n398), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT81), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n290), .B1(new_n316), .B2(G33), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n297), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n222), .B1(new_n418), .B2(new_n288), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n404), .B1(new_n419), .B2(new_n402), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n261), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT81), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n398), .ZN(new_n423));
  MUX2_X1   g0223(.A(G223), .B(G226), .S(G1698), .Z(new_n424));
  NAND2_X1  g0224(.A1(new_n317), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n338), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n336), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n375), .B2(new_n339), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n336), .B1(G232), .B2(new_n340), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n317), .A2(new_n424), .B1(G33), .B2(G87), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(G179), .C1(new_n338), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n414), .A2(new_n423), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n427), .B2(new_n429), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n431), .B(G190), .C1(new_n338), .C2(new_n432), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(new_n421), .A3(new_n398), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n299), .A2(G68), .ZN(new_n443));
  INV_X1    g0243(.A(new_n402), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n262), .B1(new_n445), .B2(new_n404), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n397), .B1(new_n446), .B2(new_n416), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT17), .A3(new_n439), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n436), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT13), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n339), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(G238), .B1(new_n339), .B2(new_n454), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n428), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n314), .A2(new_n290), .A3(G226), .A4(new_n309), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n314), .A2(new_n290), .A3(G232), .A4(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G97), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n460), .A2(new_n461), .A3(new_n465), .A4(new_n462), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n453), .B(new_n459), .C1(new_n467), .C2(new_n338), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n338), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT13), .B1(new_n469), .B2(new_n458), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(G179), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n472), .A3(new_n470), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n469), .A2(new_n458), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT77), .A3(new_n453), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(G169), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT14), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n473), .A2(KEYINPUT14), .A3(G169), .A4(new_n475), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n382), .A2(new_n202), .B1(new_n212), .B2(G68), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n385), .A2(new_n227), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n261), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT11), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT12), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n356), .B2(new_n222), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n358), .A2(new_n222), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR3_X1    g0290(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n480), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n473), .A2(G200), .A3(new_n475), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n393), .B1(new_n474), .B2(new_n453), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n495), .B2(new_n470), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n494), .B2(new_n496), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR4_X1   g0300(.A1(new_n395), .A2(new_n452), .A3(new_n493), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n307), .A2(KEYINPUT86), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT86), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n269), .C1(new_n305), .C2(new_n306), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n329), .A2(new_n346), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G190), .B2(new_n329), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n338), .A2(new_n211), .A3(G45), .A4(G274), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n338), .A2(G250), .A3(new_n321), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT87), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT87), .B1(new_n508), .B2(new_n509), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G238), .A2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n228), .B2(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n408), .A3(new_n314), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT88), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G33), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n338), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n512), .A2(new_n393), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n522), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n346), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n384), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n263), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n265), .A2(new_n224), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n408), .A2(new_n212), .A3(G68), .A4(new_n314), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n212), .B1(new_n462), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n272), .A2(new_n224), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n537), .A2(new_n538), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT89), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n262), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(KEYINPUT89), .A3(new_n540), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n533), .B(new_n534), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n266), .A2(new_n532), .ZN(new_n546));
  INV_X1    g0346(.A(new_n533), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n512), .B2(new_n522), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n528), .A2(new_n529), .A3(G179), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n531), .A2(new_n544), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT93), .ZN(new_n553));
  XOR2_X1   g0353(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n554));
  NOR2_X1   g0354(.A1(new_n263), .A2(G107), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n206), .B2(new_n265), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n206), .A2(G20), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n520), .A2(new_n212), .A3(G33), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n224), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n317), .A2(new_n212), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n212), .A2(G87), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n564), .B1(new_n374), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n560), .A3(new_n561), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n212), .A2(new_n408), .A3(new_n314), .A4(new_n565), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT24), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n557), .B1(new_n573), .B2(new_n261), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n325), .A2(G264), .B1(new_n327), .B2(new_n324), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n217), .B2(G1698), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n408), .A3(new_n314), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G294), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n575), .B(new_n331), .C1(new_n580), .C2(new_n338), .ZN(new_n581));
  INV_X1    g0381(.A(new_n324), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G264), .A3(new_n338), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n327), .A2(new_n324), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n338), .B1(new_n578), .B2(new_n579), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n380), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n553), .B1(new_n574), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n581), .A2(new_n587), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n262), .B1(new_n569), .B2(new_n572), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(KEYINPUT93), .C1(new_n591), .C2(new_n557), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n585), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G190), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n585), .B2(new_n586), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n574), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n552), .A2(new_n589), .A3(new_n592), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n325), .A2(G270), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n584), .ZN(new_n599));
  NOR2_X1   g0399(.A1(G257), .A2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n218), .B2(G1698), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n408), .A3(new_n314), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n374), .A2(G303), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n308), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(KEYINPUT90), .A3(new_n308), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n599), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n311), .B(new_n212), .C1(G33), .C2(new_n205), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n261), .B(new_n610), .C1(new_n520), .C2(new_n212), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT20), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n265), .A2(new_n516), .B1(new_n520), .B2(new_n263), .ZN(new_n613));
  OAI21_X1  g0413(.A(G169), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT21), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n599), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT90), .B1(new_n604), .B2(new_n308), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n606), .B(new_n338), .C1(new_n602), .C2(new_n603), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(new_n613), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n611), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(new_n620), .A3(G169), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G179), .B1(new_n612), .B2(new_n613), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT91), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n331), .B1(new_n621), .B2(new_n623), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n609), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n619), .B2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n609), .A2(G190), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n626), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n597), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n333), .A2(new_n501), .A3(new_n507), .A4(new_n637), .ZN(G372));
  AND2_X1   g0438(.A1(new_n494), .A2(new_n496), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n390), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n450), .B1(new_n493), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n434), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n421), .B2(new_n398), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n367), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n370), .ZN(new_n647));
  INV_X1    g0447(.A(new_n548), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n596), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n531), .A2(new_n544), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n626), .A2(new_n632), .ZN(new_n655));
  INV_X1    g0455(.A(new_n574), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n590), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n654), .A2(new_n658), .A3(new_n507), .A4(new_n333), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n307), .A2(new_n332), .A3(new_n552), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n651), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n651), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n502), .A2(new_n504), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n332), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n659), .B(new_n661), .C1(KEYINPUT26), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n501), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n647), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n624), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n655), .A2(new_n635), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n655), .B2(new_n674), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT95), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT95), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n589), .A2(new_n592), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n596), .ZN(new_n684));
  INV_X1    g0484(.A(new_n673), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n574), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n657), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n655), .A2(new_n673), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n657), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n685), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n216), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n538), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n233), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n655), .A2(new_n683), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n654), .A2(new_n702), .A3(new_n507), .A4(new_n333), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n551), .B(KEYINPUT94), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n548), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n307), .A2(new_n552), .A3(new_n707), .A4(new_n332), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n651), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n701), .A2(new_n703), .A3(new_n712), .ZN(new_n713));
  AND4_X1   g0513(.A1(KEYINPUT97), .A2(new_n713), .A3(KEYINPUT29), .A4(new_n685), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n673), .B1(new_n715), .B2(new_n703), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT97), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n665), .A2(new_n685), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n714), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n637), .A2(new_n507), .A3(new_n333), .A4(new_n685), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n329), .A2(new_n550), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n607), .A2(new_n608), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n593), .A2(new_n598), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n512), .A2(new_n522), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(G179), .A3(new_n320), .A4(new_n328), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n593), .B(new_n598), .C1(new_n617), .C2(new_n618), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n729), .A2(new_n593), .A3(G179), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n329), .A3(new_n619), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n673), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n722), .B1(new_n723), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n721), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n700), .B1(new_n741), .B2(new_n211), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(G364));
  AND2_X1   g0543(.A1(new_n212), .A2(G13), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n211), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n694), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n679), .A2(new_n722), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n681), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n260), .B1(G20), .B2(new_n380), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT100), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n253), .A2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(G45), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n233), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n408), .A2(new_n314), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n215), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n760), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n216), .A2(new_n374), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n516), .B2(new_n216), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n759), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G20), .A3(new_n393), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G329), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n212), .A2(new_n331), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n393), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n287), .B(new_n779), .C1(G311), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n774), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n393), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G326), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n782), .A2(G190), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n212), .A2(new_n393), .A3(new_n346), .A4(G179), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(new_n786), .B1(G303), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n212), .B1(new_n770), .B2(G190), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n212), .A2(new_n346), .A3(G179), .A4(G190), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(G294), .B1(new_n791), .B2(G283), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n781), .A2(new_n784), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(G97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n780), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n795), .B2(new_n227), .C1(new_n250), .C2(new_n777), .ZN(new_n796));
  INV_X1    g0596(.A(new_n783), .ZN(new_n797));
  INV_X1    g0597(.A(new_n785), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n202), .A2(new_n797), .B1(new_n798), .B2(new_n222), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n206), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n772), .A2(G159), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(KEYINPUT32), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n800), .B(new_n804), .C1(KEYINPUT32), .C2(new_n803), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n787), .A2(G87), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n287), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT101), .Z(new_n808));
  OAI21_X1  g0608(.A(new_n793), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n769), .B(new_n748), .C1(new_n809), .C2(new_n754), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n757), .B(KEYINPUT102), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n680), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n750), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT103), .Z(G396));
  NAND2_X1  g0614(.A1(new_n389), .A2(new_n673), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n394), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n390), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n390), .A2(new_n673), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n718), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n665), .A2(new_n685), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n747), .B1(new_n823), .B2(new_n740), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n740), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n754), .A2(new_n755), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n747), .B1(new_n827), .B2(G77), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n777), .A2(new_n829), .B1(new_n830), .B2(new_n771), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n287), .B(new_n831), .C1(new_n520), .C2(new_n780), .ZN(new_n832));
  INV_X1    g0632(.A(G303), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT104), .B(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n833), .A2(new_n797), .B1(new_n798), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G107), .B2(new_n787), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n791), .A2(G87), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n832), .A2(new_n794), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G143), .A2(new_n776), .B1(new_n780), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n797), .C1(new_n841), .C2(new_n798), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n791), .A2(G68), .ZN(new_n846));
  INV_X1    g0646(.A(new_n787), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n250), .B2(new_n789), .C1(new_n847), .C2(new_n202), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n763), .B(new_n848), .C1(G132), .C2(new_n772), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n838), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n828), .B1(new_n851), .B2(new_n754), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n821), .B2(new_n756), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n825), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  INV_X1    g0655(.A(KEYINPUT107), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n763), .A2(new_n286), .A3(new_n212), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n411), .A2(G68), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n405), .B1(new_n858), .B2(new_n444), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n262), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT107), .B(new_n261), .C1(new_n415), .C2(new_n405), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n416), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n642), .B1(new_n862), .B2(new_n398), .ZN(new_n863));
  INV_X1    g0663(.A(new_n440), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT108), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT108), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n261), .B1(new_n415), .B2(new_n405), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n412), .B1(new_n867), .B2(new_n856), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n397), .B1(new_n868), .B2(new_n861), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n866), .B(new_n440), .C1(new_n869), .C2(new_n642), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n671), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n671), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n414), .A2(new_n423), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n447), .B2(new_n439), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n435), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT109), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n435), .A2(new_n874), .A3(KEYINPUT109), .A4(new_n875), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n872), .A2(KEYINPUT37), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n449), .B1(KEYINPUT18), .B2(new_n435), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n871), .B1(new_n882), .B2(new_n436), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n864), .A2(new_n643), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n874), .B1(new_n644), .B2(new_n450), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n881), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT110), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT110), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n881), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n884), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n480), .B1(new_n499), .B2(new_n498), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n492), .A2(new_n685), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n639), .A2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n480), .B2(new_n492), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n819), .B1(new_n723), .B2(new_n738), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n881), .B1(new_n880), .B2(new_n883), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n869), .A2(new_n671), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n452), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n440), .B1(new_n869), .B2(new_n642), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(KEYINPUT108), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n885), .B1(new_n908), .B2(new_n870), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n878), .A2(new_n879), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT38), .B(new_n906), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n903), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n894), .A2(new_n902), .B1(new_n912), .B2(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n723), .A2(new_n738), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n501), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n722), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT111), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n913), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n647), .ZN(new_n922));
  INV_X1    g0722(.A(new_n721), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n501), .ZN(new_n924));
  INV_X1    g0724(.A(new_n493), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n673), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n904), .A2(new_n911), .A3(KEYINPUT39), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n894), .C2(KEYINPUT39), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n644), .A2(new_n873), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n897), .A2(new_n899), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n822), .B2(new_n818), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n904), .A2(new_n911), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n924), .B(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n921), .A2(new_n935), .B1(new_n211), .B2(new_n744), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n921), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n233), .B(G77), .C1(new_n250), .C2(new_n222), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n202), .A2(G68), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n211), .B(G13), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n260), .A2(new_n212), .A3(new_n516), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n279), .A2(new_n284), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT105), .Z(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT35), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  XNOR2_X1  g0747(.A(KEYINPUT106), .B(KEYINPUT36), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n937), .A2(new_n940), .A3(new_n949), .ZN(G367));
  INV_X1    g0750(.A(G159), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n798), .A2(new_n951), .B1(new_n250), .B2(new_n847), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G68), .B2(new_n790), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n374), .B1(new_n772), .B2(G137), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G50), .A2(new_n780), .B1(new_n776), .B2(G150), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n783), .A2(G143), .B1(G77), .B2(new_n791), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n795), .A2(new_n834), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n317), .B(new_n958), .C1(G317), .C2(new_n772), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT46), .B1(new_n847), .B2(new_n516), .ZN(new_n960));
  INV_X1    g0760(.A(new_n520), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n962), .B2(new_n847), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n798), .A2(new_n829), .B1(new_n205), .B2(new_n801), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G107), .B2(new_n790), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n959), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n776), .A2(G303), .B1(new_n783), .B2(G311), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT112), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n957), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT47), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n754), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n765), .A2(new_n247), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n758), .B1(new_n215), .B2(new_n384), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n747), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT113), .Z(new_n977));
  OR2_X1    g0777(.A1(new_n544), .A2(new_n685), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n662), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n705), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n811), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n694), .B(KEYINPUT41), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n663), .A2(new_n673), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n333), .A3(new_n507), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n663), .A2(new_n332), .A3(new_n673), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n692), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n692), .A2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n682), .A3(new_n687), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n688), .A3(new_n990), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n690), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n687), .B2(new_n689), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n681), .B(new_n996), .Z(new_n997));
  INV_X1    g0797(.A(new_n741), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n994), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n982), .B1(new_n1001), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n746), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n986), .A2(new_n690), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT42), .Z(new_n1005));
  INV_X1    g0805(.A(new_n986), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n333), .B1(new_n1006), .B2(new_n683), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n685), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1005), .A2(new_n1008), .B1(KEYINPUT43), .B2(new_n980), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n688), .A2(new_n1006), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n981), .B1(new_n1003), .B2(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(new_n696), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n767), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(G107), .B2(new_n215), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n244), .A2(G45), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n765), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n351), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  AOI211_X1 g0821(.A(G45), .B(new_n1015), .C1(G68), .C2(G77), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1017), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n747), .B1(new_n1024), .B2(new_n759), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n847), .A2(new_n829), .B1(new_n789), .B2(new_n834), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G303), .A2(new_n780), .B1(new_n776), .B2(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n830), .B2(new_n798), .C1(new_n778), .C2(new_n797), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n801), .A2(new_n961), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n317), .B(new_n1035), .C1(G326), .C2(new_n772), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n317), .B1(new_n841), .B2(new_n771), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n847), .A2(new_n227), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G97), .C2(new_n791), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT114), .Z(new_n1041));
  NOR2_X1   g0841(.A1(new_n789), .A2(new_n384), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n776), .B2(G50), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT115), .Z(new_n1044));
  OAI22_X1  g0844(.A1(new_n795), .A2(new_n222), .B1(new_n797), .B2(new_n951), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n352), .B2(new_n785), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1041), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1025), .B1(new_n1048), .B2(new_n754), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n687), .B2(new_n811), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT116), .Z(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n997), .B2(new_n746), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n999), .A2(new_n694), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n997), .A2(new_n998), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  AOI21_X1  g0855(.A(new_n695), .B1(new_n994), .B2(new_n1000), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1000), .B2(new_n994), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n994), .A2(new_n746), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n754), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n776), .A2(G159), .B1(new_n783), .B2(G150), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT51), .Z(new_n1061));
  NOR2_X1   g0861(.A1(new_n795), .A2(new_n351), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n763), .B(new_n1062), .C1(G143), .C2(new_n772), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n789), .A2(new_n227), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n837), .B1(new_n847), .B2(new_n222), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G50), .C2(new_n785), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1061), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n776), .A2(G311), .B1(new_n783), .B2(G317), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n374), .B1(new_n771), .B2(new_n778), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n780), .B2(G294), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n798), .A2(new_n833), .B1(new_n789), .B2(new_n961), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n847), .A2(new_n834), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n802), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1059), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n758), .B1(new_n205), .B2(new_n215), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n257), .B2(new_n765), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n748), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n757), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n986), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1057), .A2(new_n1058), .A3(new_n1081), .ZN(G390));
  NAND2_X1  g0882(.A1(new_n891), .A2(new_n893), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n911), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n926), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n818), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n716), .B2(new_n817), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1085), .C1(new_n930), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n927), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT39), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n931), .A2(new_n926), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n900), .A2(new_n901), .A3(G330), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1088), .B(new_n1094), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n746), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n747), .B1(new_n827), .B2(new_n352), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n795), .A2(new_n205), .B1(new_n771), .B2(new_n829), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n287), .B(new_n1100), .C1(G116), .C2(new_n776), .ZN(new_n1101));
  INV_X1    g0901(.A(G283), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n797), .A2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1064), .B(new_n1103), .C1(G107), .C2(new_n785), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1104), .A3(new_n806), .A4(new_n846), .ZN(new_n1105));
  INV_X1    g0905(.A(G132), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1106), .A2(new_n777), .B1(new_n795), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n374), .B(new_n1108), .C1(G125), .C2(new_n772), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n785), .A2(G137), .B1(G50), .B2(new_n791), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n783), .A2(G128), .B1(G159), .B2(new_n790), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n787), .A2(G150), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1105), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1115), .B2(new_n754), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT119), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1091), .B2(new_n756), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1098), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1098), .A2(new_n1121), .A3(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n501), .A2(new_n739), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n501), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n647), .B(new_n1125), .C1(new_n721), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n722), .B(new_n819), .C1(new_n723), .C2(new_n738), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n900), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n901), .A2(G330), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(KEYINPUT117), .A3(new_n930), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1087), .A2(new_n1130), .A3(new_n1094), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n713), .A2(new_n685), .A3(new_n817), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1094), .A2(new_n1135), .A3(new_n818), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT118), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n822), .A2(new_n818), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1129), .A2(new_n900), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1095), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1127), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n695), .B1(new_n1124), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1096), .A2(new_n1143), .A3(new_n1097), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1147), .ZN(G378));
  OR2_X1    g0948(.A1(new_n317), .A2(G41), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n795), .A2(new_n384), .B1(new_n771), .B2(new_n1102), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G107), .C2(new_n776), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n783), .A2(G116), .B1(G68), .B2(new_n790), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT121), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n801), .A2(new_n250), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1154), .B(new_n1039), .C1(G97), .C2(new_n785), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT58), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1149), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n783), .A2(G125), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n798), .B2(new_n1106), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G128), .A2(new_n776), .B1(new_n780), .B2(G137), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n847), .B2(new_n1107), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n790), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n791), .A2(G159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1160), .B1(KEYINPUT58), .B2(new_n1157), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1172), .A2(new_n754), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n747), .B1(new_n827), .B2(G50), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n370), .B1(new_n365), .B2(new_n366), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n360), .A2(new_n671), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1178), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n367), .A2(new_n370), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n1179), .A3(new_n1175), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1182), .A2(KEYINPUT122), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT122), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1173), .B(new_n1174), .C1(new_n1188), .C2(new_n755), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1190));
  OAI21_X1  g0990(.A(G330), .B1(new_n894), .B2(new_n902), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n912), .A2(KEYINPUT40), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT123), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT123), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1195), .B(new_n1190), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1191), .A2(new_n1192), .A3(new_n1188), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n934), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1198), .A2(new_n934), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1197), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT124), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1189), .B1(new_n1205), .B2(new_n746), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1127), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1146), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT57), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1200), .A2(new_n934), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n694), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1209), .B2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n746), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n748), .B1(new_n826), .B2(new_n222), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n287), .B1(new_n772), .B2(G303), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n795), .B2(new_n206), .C1(new_n1102), .C2(new_n777), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1042), .B(new_n1218), .C1(G77), .C2(new_n791), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n829), .A2(new_n797), .B1(new_n798), .B2(new_n961), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G97), .B2(new_n787), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n780), .A2(G150), .B1(G128), .B2(new_n772), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n840), .B2(new_n777), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1223), .A2(new_n763), .A3(new_n1154), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n797), .A2(new_n1106), .B1(new_n951), .B2(new_n847), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n798), .A2(new_n1107), .B1(new_n202), .B2(new_n789), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1219), .A2(new_n1221), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1216), .B1(new_n1059), .B2(new_n1228), .C1(new_n900), .C2(new_n756), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1215), .A2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n982), .B(KEYINPUT125), .Z(new_n1231));
  NOR2_X1   g1031(.A1(new_n1143), .A2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1127), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(G381));
  NOR2_X1   g1036(.A1(G387), .A2(G390), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OR3_X1    g1038(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1235), .A3(new_n1241), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G378), .A2(new_n1238), .A3(new_n1242), .A4(G375), .ZN(G407));
  AOI22_X1  g1043(.A1(new_n1120), .A2(new_n1122), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n672), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  AOI21_X1  g1048(.A(KEYINPUT60), .B1(new_n1233), .B2(new_n1127), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(new_n695), .A3(new_n1143), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1139), .A2(new_n1127), .A3(KEYINPUT60), .A4(new_n1142), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1251), .B(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1230), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n854), .B(new_n1230), .C1(new_n1250), .C2(new_n1253), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G2897), .B(new_n1246), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n854), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1254), .A2(G384), .A3(new_n1255), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1246), .A2(G2897), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1206), .C1(new_n1209), .C2(new_n1212), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n934), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1196), .ZN(new_n1269));
  OAI221_X1 g1069(.A(G330), .B1(new_n912), .B2(KEYINPUT40), .C1(new_n894), .C2(new_n902), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1195), .B1(new_n1270), .B2(new_n1190), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1202), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1197), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1268), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1208), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1231), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1189), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1211), .B2(new_n745), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1244), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1266), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1245), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(G393), .B(G396), .Z(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(G390), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1292), .B2(new_n1237), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1238), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1246), .B1(new_n1266), .B2(new_n1281), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1286), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1284), .A2(new_n1288), .A3(new_n1295), .A4(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1296), .A2(new_n1299), .A3(new_n1286), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1296), .B2(new_n1264), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1296), .B2(new_n1286), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1298), .B1(new_n1304), .B2(new_n1295), .ZN(G405));
  AND2_X1   g1105(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G375), .A2(new_n1244), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1266), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1286), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1287), .A3(new_n1266), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1306), .B(new_n1311), .ZN(G402));
endmodule


