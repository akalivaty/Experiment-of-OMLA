//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT18), .A3(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT18), .A2(G131), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n193), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G125), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(new_n197), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT84), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n195), .A2(new_n207), .A3(new_n197), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G113), .B(G122), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT16), .ZN(new_n216));
  OR3_X1    g030(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G146), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(G146), .B1(new_n216), .B2(new_n217), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n194), .A2(KEYINPUT17), .A3(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n194), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n191), .A2(new_n224), .A3(new_n193), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n221), .B(new_n222), .C1(new_n226), .C2(KEYINPUT17), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n212), .A2(new_n215), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n202), .A2(KEYINPUT19), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT19), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n204), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n232), .A3(new_n205), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n229), .A2(new_n235), .B1(new_n209), .B2(new_n211), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n236), .B2(new_n215), .ZN(new_n237));
  NOR2_X1   g051(.A1(G475), .A2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT20), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT87), .B1(new_n190), .B2(G128), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n190), .A2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT88), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT13), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n190), .A2(KEYINPUT13), .A3(G128), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G134), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G122), .ZN(new_n259));
  INV_X1    g073(.A(G122), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G116), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G107), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G107), .B1(new_n259), .B2(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT88), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n248), .A2(new_n267), .A3(new_n249), .A4(new_n250), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n252), .A2(new_n257), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n258), .A2(G122), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n259), .B1(KEYINPUT14), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n270), .A2(KEYINPUT14), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n271), .B2(new_n272), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n263), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n251), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n249), .B1(new_n248), .B2(new_n250), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n264), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n269), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT9), .B(G234), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(G217), .A3(new_n188), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  INV_X1    g099(.A(new_n283), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n269), .B(new_n286), .C1(new_n276), .C2(new_n279), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n280), .A2(KEYINPUT90), .A3(new_n283), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G478), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT15), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n291), .A2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(new_n228), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n215), .B1(new_n212), .B2(new_n227), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT86), .B(G475), .Z(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n243), .A2(new_n294), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n188), .A2(G952), .ZN(new_n302));
  INV_X1    g116(.A(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(new_n187), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(G902), .B(G953), .C1(new_n303), .C2(new_n187), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT91), .Z(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT21), .B(G898), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT92), .B1(new_n301), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n295), .A2(new_n294), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n240), .A2(new_n242), .B1(new_n298), .B2(new_n299), .ZN(new_n313));
  INV_X1    g127(.A(new_n309), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT2), .B(G113), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT66), .A2(G119), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n258), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n322), .A2(G116), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT67), .B1(new_n325), .B2(new_n326), .ZN(new_n328));
  AND2_X1   g142(.A1(KEYINPUT66), .A2(G119), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT66), .A2(G119), .ZN(new_n330));
  OAI21_X1  g144(.A(G116), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n332));
  INV_X1    g146(.A(new_n326), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G113), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n325), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n327), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n214), .A2(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n263), .A2(G104), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT77), .B1(new_n263), .B2(G104), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n214), .A3(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n263), .A3(G104), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n340), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT78), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n348), .A2(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n340), .A4(new_n347), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n343), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n339), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT81), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n339), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G101), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n352), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n340), .B1(new_n353), .B2(new_n347), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(KEYINPUT79), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n325), .A2(KEYINPUT67), .A3(new_n326), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n320), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n325), .A2(new_n326), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n319), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n364), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n358), .A2(new_n360), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(G110), .B(G122), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n358), .A2(new_n379), .A3(new_n375), .A4(new_n360), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n382), .A3(new_n377), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n205), .A2(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n190), .A2(G146), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT0), .A4(G128), .ZN(new_n386));
  XNOR2_X1  g200(.A(G143), .B(G146), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G128), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G125), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(new_n246), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT64), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(new_n387), .B2(new_n396), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n395), .A2(new_n396), .A3(new_n384), .A4(new_n385), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n390), .B1(new_n399), .B2(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n188), .A2(G224), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND3_X1  g216(.A1(new_n381), .A2(new_n383), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(KEYINPUT7), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n380), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n377), .B(KEYINPUT8), .Z(new_n410));
  NOR2_X1   g224(.A1(new_n339), .A2(new_n356), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n327), .B1(new_n413), .B2(new_n338), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n356), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n411), .B2(KEYINPUT82), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n410), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n403), .A2(new_n420), .A3(new_n418), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n318), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G221), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n282), .B2(new_n289), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n426), .B(KEYINPUT76), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n289), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  INV_X1    g245(.A(G227), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n431), .B(new_n433), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n352), .A2(new_n355), .ZN(new_n436));
  INV_X1    g250(.A(new_n343), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n392), .A2(KEYINPUT80), .ZN(new_n438));
  OAI21_X1  g252(.A(G128), .B1(new_n392), .B2(KEYINPUT80), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n391), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n396), .A2(new_n384), .A3(new_n385), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT64), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n387), .A2(new_n395), .A3(new_n396), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n436), .A2(new_n437), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n392), .A2(G128), .B1(new_n384), .B2(new_n385), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n442), .B2(new_n443), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n447), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n446), .A2(new_n447), .B1(new_n450), .B2(new_n356), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT11), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n249), .B2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT11), .A3(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n249), .A2(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(new_n224), .A4(new_n456), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n389), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n367), .A2(new_n461), .A3(new_n374), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n451), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n451), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n435), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n436), .A2(new_n437), .A3(new_n445), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n399), .B1(new_n436), .B2(new_n437), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT12), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n451), .A2(new_n460), .A3(new_n462), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n434), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n430), .B1(new_n475), .B2(new_n429), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n435), .ZN(new_n478));
  INV_X1    g292(.A(new_n464), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n471), .A3(new_n434), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n480), .A3(G469), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n428), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n316), .A2(new_n424), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(G472), .A2(G902), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n249), .A2(G137), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n454), .A2(G134), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n459), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n399), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n461), .A2(new_n466), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n372), .A3(new_n493), .A4(new_n370), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n449), .B2(new_n490), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n399), .A2(KEYINPUT65), .A3(new_n491), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n493), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n373), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n494), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n497), .B1(new_n503), .B2(KEYINPUT28), .ZN(new_n504));
  AOI211_X1 g318(.A(KEYINPUT69), .B(new_n495), .C1(new_n502), .C2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n192), .A2(G210), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(G101), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n490), .B1(new_n444), .B2(new_n394), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n389), .B1(new_n458), .B2(new_n459), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n516), .A3(new_n373), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n494), .A2(new_n509), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n515), .B1(new_n511), .B2(new_n501), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n518), .B1(new_n523), .B2(new_n373), .ZN(new_n524));
  NOR2_X1   g338(.A1(KEYINPUT68), .A2(KEYINPUT31), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n486), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT69), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n319), .B1(new_n328), .B2(new_n334), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n327), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n514), .B1(new_n492), .B2(new_n498), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n500), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n460), .A2(new_n389), .B1(new_n449), .B2(new_n490), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n373), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n530), .B(KEYINPUT28), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n509), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n495), .B1(new_n502), .B2(new_n494), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n497), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n525), .B1(new_n517), .B2(new_n519), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n522), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n544));
  OAI22_X1  g358(.A1(new_n513), .A2(new_n514), .B1(new_n531), .B2(new_n327), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n494), .A2(new_n545), .A3(KEYINPUT71), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n373), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(KEYINPUT28), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n538), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n496), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n552), .A2(new_n289), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n530), .B1(new_n494), .B2(new_n495), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n536), .B1(new_n373), .B2(new_n501), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n495), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n538), .B1(new_n556), .B2(new_n537), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n536), .B1(new_n523), .B2(new_n373), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n550), .B1(new_n558), .B2(new_n509), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n553), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n529), .A2(new_n544), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G217), .B1(new_n303), .B2(G902), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT72), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n323), .A2(new_n246), .A3(new_n324), .ZN(new_n566));
  AND2_X1   g380(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n567));
  NOR2_X1   g381(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n246), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT73), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n246), .A3(KEYINPUT23), .A4(G119), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G110), .ZN(new_n576));
  OAI21_X1  g390(.A(G128), .B1(new_n329), .B2(new_n330), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n246), .B1(new_n323), .B2(new_n324), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n566), .B2(new_n569), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n576), .A4(new_n575), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  NAND2_X1  g398(.A1(new_n246), .A2(G119), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n577), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n218), .A2(new_n206), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n577), .A2(new_n585), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n219), .B2(new_n220), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n576), .B1(new_n581), .B2(new_n575), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT22), .B(G137), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n425), .A2(new_n303), .A3(G953), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n586), .B1(new_n578), .B2(KEYINPUT75), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n589), .B1(new_n602), .B2(new_n583), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n594), .A2(new_n595), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n289), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n601), .A2(new_n605), .A3(KEYINPUT25), .A4(new_n289), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n565), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n601), .A2(new_n605), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n303), .B2(G217), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n562), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n483), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n340), .ZN(G3));
  AOI211_X1 g431(.A(new_n518), .B(new_n520), .C1(new_n523), .C2(new_n373), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n541), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n619), .B2(new_n540), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n527), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n614), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n482), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT93), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n237), .A2(new_n241), .A3(new_n238), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n241), .B1(new_n237), .B2(new_n238), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n300), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n291), .A2(new_n292), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n288), .A2(new_n631), .A3(new_n290), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n284), .A2(KEYINPUT33), .A3(new_n287), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n289), .A2(G478), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n629), .A2(new_n636), .A3(new_n314), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n403), .A2(new_n420), .A3(new_n418), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n420), .B1(new_n403), .B2(new_n418), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n637), .B(new_n317), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  XNOR2_X1  g458(.A(new_n309), .B(KEYINPUT94), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n317), .B(new_n645), .C1(new_n638), .C2(new_n639), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n311), .A2(new_n629), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n608), .A2(new_n609), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n564), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n591), .A2(new_n596), .A3(new_n656), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n603), .A2(new_n604), .B1(KEYINPUT36), .B2(new_n599), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n613), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n653), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n660), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n610), .A2(new_n662), .A3(KEYINPUT95), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n622), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n316), .A3(new_n424), .A4(new_n482), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NOR2_X1   g481(.A1(new_n661), .A2(new_n663), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n424), .A2(new_n562), .A3(new_n482), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n305), .B1(new_n307), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n648), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n246), .ZN(G30));
  AOI211_X1 g489(.A(new_n528), .B(new_n485), .C1(new_n619), .C2(new_n540), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT32), .B1(new_n543), .B2(new_n486), .ZN(new_n677));
  INV_X1    g491(.A(new_n558), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n509), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n546), .A2(new_n548), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(new_n538), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n621), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n676), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n311), .A2(new_n313), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n683), .A2(new_n668), .A3(new_n684), .A4(new_n318), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n638), .A2(new_n639), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n422), .A2(new_n423), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT38), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n671), .B(KEYINPUT39), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n482), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n685), .A2(new_n692), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND2_X1  g513(.A1(new_n629), .A2(new_n636), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n671), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n669), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n205), .ZN(G48));
  NOR2_X1   g518(.A1(new_n676), .A2(new_n677), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n623), .B1(new_n705), .B2(new_n561), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n465), .A2(new_n474), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n289), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n429), .A3(new_n289), .ZN(new_n710));
  INV_X1    g524(.A(new_n426), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n706), .A2(new_n641), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT96), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  OAI21_X1  g531(.A(new_n317), .B1(new_n638), .B2(new_n639), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n712), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n649), .A2(new_n706), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n562), .A3(new_n316), .A4(new_n668), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  INV_X1    g537(.A(new_n646), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n712), .A2(new_n684), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n549), .A2(new_n496), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n538), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n485), .B1(new_n619), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT97), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n620), .B2(new_n621), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n289), .B1(new_n510), .B2(new_n526), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT97), .A3(G472), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n724), .A2(new_n725), .A3(new_n733), .A4(new_n614), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n732), .ZN(new_n736));
  INV_X1    g550(.A(new_n728), .ZN(new_n737));
  AND4_X1   g551(.A1(KEYINPUT98), .A2(new_n736), .A3(new_n668), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT98), .B1(new_n733), .B2(new_n668), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n701), .B(new_n719), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND2_X1  g555(.A1(new_n478), .A2(new_n480), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n463), .A2(new_n464), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT99), .B1(new_n744), .B2(new_n434), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(G469), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n426), .B1(new_n747), .B2(new_n476), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n638), .A2(new_n639), .A3(new_n318), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n706), .A2(new_n701), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT42), .B1(new_n750), .B2(KEYINPUT100), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n224), .ZN(G33));
  NAND3_X1  g569(.A1(new_n706), .A2(new_n748), .A3(new_n749), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n673), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n249), .ZN(G36));
  NAND2_X1  g572(.A1(new_n686), .A2(new_n317), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n313), .A2(new_n636), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT43), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n622), .A3(new_n668), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n743), .A2(KEYINPUT45), .A3(new_n746), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n429), .B1(new_n742), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n430), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n771), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT101), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .B1(new_n429), .B2(new_n475), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n711), .A3(new_n694), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT102), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(KEYINPUT102), .A3(new_n711), .A4(new_n694), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n767), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n454), .ZN(G39));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n711), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n775), .A2(new_n784), .A3(new_n711), .ZN(new_n785));
  INV_X1    g599(.A(new_n671), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n749), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n562), .A2(new_n614), .A3(new_n700), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n783), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n198), .ZN(G42));
  XNOR2_X1  g605(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n691), .A2(new_n318), .A3(new_n713), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n733), .A2(new_n614), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n304), .B1(new_n761), .B2(new_n762), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n794), .A2(new_n795), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n793), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n805), .B(new_n793), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n802), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n800), .A3(KEYINPUT50), .A4(new_n796), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n801), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT116), .A3(KEYINPUT50), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n807), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n759), .A2(new_n712), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n614), .A3(new_n305), .A4(new_n683), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n629), .A3(new_n636), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n798), .A2(new_n817), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT97), .B1(new_n731), .B2(G472), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n729), .B(new_n621), .C1(new_n543), .C2(new_n289), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n668), .B(new_n737), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT98), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n733), .A2(KEYINPUT98), .A3(new_n668), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n819), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n709), .A2(new_n710), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n427), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT113), .Z(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n783), .B2(new_n785), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n799), .A2(new_n759), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n792), .B1(new_n816), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n820), .A2(new_n706), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  INV_X1    g655(.A(new_n719), .ZN(new_n842));
  OAI221_X1 g656(.A(new_n302), .B1(new_n799), .B2(new_n842), .C1(new_n700), .C2(new_n818), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n833), .B1(new_n783), .B2(new_n785), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n836), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT51), .B(new_n831), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(new_n807), .B2(new_n814), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(new_n753), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n720), .A2(new_n722), .A3(new_n714), .A4(new_n734), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n751), .ZN(new_n858));
  INV_X1    g672(.A(new_n700), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n624), .A2(new_n482), .A3(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n483), .A2(new_n615), .B1(new_n860), .B2(new_n646), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n649), .A2(new_n482), .A3(new_n624), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT104), .B1(new_n862), .B2(new_n665), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(KEYINPUT104), .A3(new_n665), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n748), .A2(new_n749), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n615), .ZN(new_n868));
  INV_X1    g682(.A(new_n301), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n562), .A2(new_n482), .A3(new_n869), .A4(new_n668), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n868), .A2(new_n672), .B1(new_n870), .B2(new_n788), .ZN(new_n871));
  INV_X1    g685(.A(new_n867), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n701), .B(new_n872), .C1(new_n738), .C2(new_n739), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT105), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n871), .B2(new_n873), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n858), .B(new_n866), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n669), .B1(new_n673), .B2(new_n702), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n702), .B1(new_n825), .B2(new_n826), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n719), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT99), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n478), .B2(new_n480), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n883), .A2(new_n429), .A3(new_n745), .ZN(new_n884));
  INV_X1    g698(.A(new_n430), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n710), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n711), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n683), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT107), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n311), .A2(new_n313), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n317), .C1(new_n638), .C2(new_n639), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n655), .A2(new_n660), .A3(new_n786), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT106), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n655), .A2(KEYINPUT106), .A3(new_n660), .A4(new_n786), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n888), .A2(new_n889), .A3(new_n892), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n682), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n529), .A2(new_n544), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n748), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT107), .B1(new_n901), .B2(new_n891), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT52), .B1(new_n881), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n669), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n672), .B2(new_n701), .ZN(new_n906));
  AND4_X1   g720(.A1(KEYINPUT52), .A2(new_n903), .A3(new_n740), .A4(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n855), .B1(new_n878), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT110), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n911), .B(new_n855), .C1(new_n878), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT111), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n855), .B1(new_n858), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n861), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n862), .A2(KEYINPUT104), .A3(new_n665), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n863), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n871), .A2(new_n873), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT105), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(new_n875), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT111), .B1(new_n754), .B2(new_n857), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n903), .A2(new_n740), .A3(new_n906), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT52), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n881), .A2(KEYINPUT52), .A3(new_n903), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT108), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n904), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n913), .A2(new_n914), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n928), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n922), .A2(new_n935), .A3(new_n858), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT53), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n922), .A2(new_n855), .A3(new_n858), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n937), .B(KEYINPUT54), .C1(new_n932), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n938), .A2(new_n932), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(KEYINPUT109), .A3(KEYINPUT54), .A4(new_n937), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n934), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n854), .A2(new_n944), .B1(G952), .B2(G953), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n623), .A2(new_n318), .A3(new_n428), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(KEYINPUT103), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(KEYINPUT103), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n900), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n832), .A2(KEYINPUT49), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n832), .A2(KEYINPUT49), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(new_n760), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n691), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n945), .A2(new_n953), .ZN(G75));
  INV_X1    g768(.A(new_n912), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n911), .B1(new_n936), .B2(new_n855), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n933), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(G210), .A3(G902), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n381), .A2(new_n383), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n402), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n958), .B2(new_n959), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n188), .A2(G952), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G51));
  XNOR2_X1  g780(.A(new_n430), .B(KEYINPUT57), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n924), .A2(new_n932), .ZN(new_n968));
  AOI211_X1 g782(.A(KEYINPUT54), .B(new_n968), .C1(new_n910), .C2(new_n912), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n914), .B1(new_n913), .B2(new_n933), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n707), .B(KEYINPUT120), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n957), .A2(G902), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n768), .A3(new_n770), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n965), .B1(new_n973), .B2(new_n976), .ZN(G54));
  INV_X1    g791(.A(new_n237), .ZN(new_n978));
  NAND2_X1  g792(.A1(KEYINPUT58), .A2(G475), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n965), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G60));
  INV_X1    g798(.A(new_n634), .ZN(new_n985));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT59), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n944), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n957), .A2(KEYINPUT54), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n934), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n989), .A2(new_n965), .A3(new_n992), .ZN(G63));
  AOI21_X1  g807(.A(new_n968), .B1(new_n910), .B2(new_n912), .ZN(new_n994));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT60), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n611), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n913), .B2(new_n933), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n965), .B1(new_n998), .B2(new_n659), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT121), .B1(new_n998), .B2(new_n659), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n997), .B(new_n999), .C1(new_n1000), .C2(KEYINPUT61), .ZN(new_n1001));
  INV_X1    g815(.A(new_n996), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n957), .A2(new_n659), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT121), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT61), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n997), .A2(new_n1003), .A3(new_n981), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1001), .A2(new_n1007), .ZN(G66));
  INV_X1    g822(.A(G224), .ZN(new_n1009));
  OAI21_X1  g823(.A(G953), .B1(new_n308), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n919), .A2(new_n857), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(G953), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n960), .B1(G898), .B2(new_n188), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(G69));
  NOR2_X1   g828(.A1(new_n188), .A2(G900), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n790), .A2(new_n780), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n778), .A2(new_n779), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(new_n706), .A3(new_n892), .ZN(new_n1018));
  INV_X1    g832(.A(new_n881), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n754), .A2(new_n1019), .A3(new_n757), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(new_n188), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n230), .A2(new_n232), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n523), .B(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT122), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n698), .A2(new_n740), .A3(new_n906), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT62), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n695), .A2(new_n759), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1029), .B(new_n706), .C1(new_n859), .C2(new_n647), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1016), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n188), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1026), .B1(new_n1032), .B2(new_n1024), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1024), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1035), .B1(new_n1031), .B2(new_n188), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n1026), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT124), .ZN(new_n1038));
  OAI21_X1  g852(.A(G953), .B1(new_n432), .B2(new_n670), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT123), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1038), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n1040), .A2(new_n1038), .ZN(new_n1043));
  OAI22_X1  g857(.A1(new_n1022), .A2(new_n1024), .B1(new_n1036), .B2(new_n1026), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1037), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1042), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1041), .A2(new_n1046), .ZN(G72));
  NAND4_X1  g861(.A1(new_n1016), .A2(new_n1011), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1048));
  NAND2_X1  g862(.A1(G472), .A2(G902), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT63), .Z(new_n1050));
  AOI21_X1  g864(.A(new_n679), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n558), .A2(new_n538), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1016), .A2(new_n1011), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1052), .B1(new_n1053), .B2(new_n1050), .ZN(new_n1054));
  NOR3_X1   g868(.A1(new_n1051), .A2(new_n1054), .A3(new_n965), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n524), .B1(new_n678), .B2(new_n538), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1050), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n942), .A2(new_n937), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT125), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n937), .A4(new_n1058), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1064), .A2(KEYINPUT126), .ZN(new_n1065));
  INV_X1    g879(.A(KEYINPUT126), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1055), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1065), .A2(new_n1067), .ZN(G57));
endmodule


