//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1103, new_n1104, new_n1105;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n459), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(G2104), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n465), .A2(KEYINPUT67), .A3(G137), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n460), .A2(new_n463), .A3(new_n466), .A4(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G2105), .B1(G101), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n472), .A2(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G112), .B2(new_n466), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n465), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND4_X1   g062(.A1(new_n466), .A2(new_n460), .A3(new_n463), .A4(new_n464), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n474), .A2(new_n464), .A3(G138), .A4(new_n466), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n460), .A2(new_n463), .A3(new_n464), .A4(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n500), .A2(KEYINPUT69), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(KEYINPUT69), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n492), .B(new_n498), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  OAI21_X1  g080(.A(G543), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(KEYINPUT70), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n509), .A2(new_n505), .A3(KEYINPUT5), .A4(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n517), .A2(G51), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n513), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n517), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n538), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT72), .B1(new_n538), .B2(new_n513), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n523), .A2(G81), .B1(G43), .B2(new_n517), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  XOR2_X1   g124(.A(KEYINPUT75), .B(G65), .Z(new_n550));
  AOI22_X1  g125(.A1(new_n511), .A2(new_n550), .B1(G78), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT76), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n513), .B1(new_n551), .B2(KEYINPUT76), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n552), .A2(new_n553), .B1(G91), .B2(new_n523), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n517), .A2(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n523), .A2(G87), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT77), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n511), .A2(G74), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n516), .A2(KEYINPUT78), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT78), .B1(new_n516), .B2(new_n565), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n564), .A2(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n523), .A2(G86), .B1(G48), .B2(new_n517), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n511), .A2(G61), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT79), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G651), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n523), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n523), .A2(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n513), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G54), .B2(new_n517), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n582), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n582), .B1(new_n589), .B2(G868), .ZN(G321));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G299), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g176(.A(G123), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n466), .A2(G111), .ZN(new_n603));
  OAI21_X1  g178(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n485), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G135), .B2(new_n488), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2096), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(G156));
  XOR2_X1   g187(.A(G1341), .B(G1348), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT81), .ZN(new_n614));
  XOR2_X1   g189(.A(G2451), .B(G2454), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT16), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n614), .B(new_n616), .Z(new_n617));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n617), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n626), .A2(G14), .A3(new_n627), .ZN(G401));
  XOR2_X1   g203(.A(G2072), .B(G2078), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT17), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2067), .B(G2678), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2084), .B(G2090), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n631), .B2(new_n632), .ZN(new_n636));
  INV_X1    g211(.A(new_n632), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(new_n633), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n634), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2096), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(G227));
  XNOR2_X1  g218(.A(G1956), .B(G2474), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1961), .B(G1966), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n644), .A3(new_n645), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n644), .B(new_n645), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n654), .B(new_n655), .C1(new_n651), .C2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1991), .B(G1996), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  INV_X1    g239(.A(G288), .ZN(new_n665));
  INV_X1    g240(.A(G16), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(G23), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT33), .B(G1976), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(G6), .A2(G16), .ZN(new_n671));
  INV_X1    g246(.A(G305), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n671), .B1(new_n672), .B2(G16), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT32), .ZN(new_n674));
  INV_X1    g249(.A(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n666), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n666), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G1971), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n668), .A2(new_n669), .ZN(new_n680));
  NAND4_X1  g255(.A1(new_n670), .A2(new_n676), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT34), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(KEYINPUT34), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n666), .A2(G24), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G290), .B2(G16), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT88), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  INV_X1    g267(.A(G119), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n466), .A2(G107), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n695));
  OAI22_X1  g270(.A1(new_n485), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G131), .B2(new_n488), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n692), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT87), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n687), .B(new_n701), .C1(new_n686), .C2(new_n685), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n682), .A2(new_n683), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT36), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n589), .A2(new_n666), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G4), .B2(new_n666), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n691), .A2(G27), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G164), .B2(new_n691), .ZN(new_n710));
  INV_X1    g285(.A(G2078), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n706), .A2(new_n707), .ZN(new_n713));
  NAND2_X1  g288(.A1(G160), .A2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G34), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT24), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n691), .B1(KEYINPUT24), .B2(new_n715), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(KEYINPUT92), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(KEYINPUT92), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n708), .A2(new_n712), .A3(new_n713), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n688), .A2(G33), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  INV_X1    g304(.A(new_n475), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n731), .B2(new_n466), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G139), .B2(new_n488), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT90), .Z(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n688), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2072), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n726), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G32), .ZN(new_n739));
  AOI21_X1  g314(.A(KEYINPUT95), .B1(new_n688), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n488), .A2(G141), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(G105), .B2(new_n478), .ZN(new_n746));
  INV_X1    g321(.A(G129), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n741), .B(new_n746), .C1(new_n747), .C2(new_n485), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n688), .ZN(new_n753));
  MUX2_X1   g328(.A(new_n740), .B(KEYINPUT95), .S(new_n753), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT96), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n666), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n666), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n606), .A2(new_n691), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT31), .B(G11), .Z(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT97), .B(G28), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(KEYINPUT30), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n764), .B2(KEYINPUT30), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G5), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G171), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1961), .ZN(new_n772));
  INV_X1    g347(.A(new_n691), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n773), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT29), .B(G2090), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(G26), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n782));
  INV_X1    g357(.A(G128), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n485), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G140), .B2(new_n488), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(new_n688), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n769), .A2(new_n772), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n666), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT23), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n543), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  NAND3_X1  g370(.A1(new_n788), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n738), .A2(new_n757), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n704), .A2(new_n798), .ZN(G311));
  INV_X1    g374(.A(G311), .ZN(G150));
  NAND2_X1  g375(.A1(new_n589), .A2(G559), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT38), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n511), .A2(G67), .ZN(new_n803));
  AND2_X1   g378(.A1(G80), .A2(G543), .ZN(new_n804));
  OAI21_X1  g379(.A(G651), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n523), .A2(G93), .B1(G55), .B2(new_n517), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(new_n542), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n802), .B(new_n811), .Z(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(G860), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  XOR2_X1   g393(.A(new_n752), .B(new_n785), .Z(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G164), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(G164), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n734), .A2(KEYINPUT100), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n734), .A2(KEYINPUT100), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n697), .B(KEYINPUT101), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n609), .ZN(new_n827));
  INV_X1    g402(.A(G130), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n466), .A2(G118), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n485), .A2(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G142), .B2(new_n488), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n823), .A2(new_n824), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n825), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n825), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n606), .B(G162), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G160), .Z(new_n839));
  AOI21_X1  g414(.A(G37), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n835), .B2(new_n836), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n844));
  OAI211_X1 g419(.A(KEYINPUT40), .B(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n842), .B(KEYINPUT102), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT40), .B1(new_n847), .B2(new_n840), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(G395));
  XOR2_X1   g424(.A(new_n588), .B(G299), .Z(new_n850));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n598), .B(new_n811), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n850), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(KEYINPUT103), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(KEYINPUT103), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n857), .A2(KEYINPUT42), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G290), .B(KEYINPUT104), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G288), .ZN(new_n861));
  XNOR2_X1  g436(.A(G303), .B(G305), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT42), .B1(new_n857), .B2(new_n858), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n859), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(G868), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n810), .A2(new_n592), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(G295));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n869), .ZN(G331));
  XNOR2_X1  g446(.A(new_n811), .B(G301), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G168), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n811), .B(G171), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G286), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n852), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n850), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n875), .B2(new_n873), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n876), .A2(new_n878), .A3(new_n863), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n863), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n884));
  NAND4_X1  g459(.A1(new_n879), .A2(new_n880), .A3(new_n884), .A4(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT44), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g465(.A(KEYINPUT106), .B(G1384), .ZN(new_n891));
  NOR2_X1   g466(.A1(G164), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT45), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n472), .A2(G40), .A3(new_n479), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n895), .A2(G1986), .A3(G290), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(G1986), .A3(G290), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT107), .ZN(new_n900));
  INV_X1    g475(.A(G1996), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n752), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n785), .B(G2067), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n697), .B(new_n700), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G1384), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT67), .B1(new_n488), .B2(G137), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n469), .A2(new_n468), .A3(new_n470), .ZN(new_n912));
  OAI211_X1 g487(.A(G40), .B(new_n479), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT69), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n500), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n497), .A2(new_n496), .ZN(new_n916));
  INV_X1    g491(.A(new_n495), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n916), .B(new_n917), .C1(new_n469), .C2(new_n490), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n908), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n910), .B1(new_n921), .B2(KEYINPUT109), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT45), .B1(new_n503), .B2(new_n908), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n913), .ZN(new_n925));
  AOI21_X1  g500(.A(G1966), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n721), .A3(new_n894), .A4(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT121), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n916), .A2(new_n917), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n469), .A2(new_n490), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n500), .B(KEYINPUT69), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n894), .B(KEYINPUT109), .C1(new_n936), .C2(KEYINPUT45), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n925), .A2(new_n937), .A3(new_n909), .ZN(new_n938));
  INV_X1    g513(.A(G1966), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT121), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n929), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n931), .A2(G8), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n931), .A2(new_n942), .A3(KEYINPUT124), .A4(G8), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(G286), .A2(G8), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT122), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT123), .B(KEYINPUT51), .Z(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n940), .B2(new_n929), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n956), .A2(KEYINPUT51), .A3(new_n949), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT126), .ZN(new_n959));
  INV_X1    g534(.A(new_n950), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n945), .B2(new_n946), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n961), .B2(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n954), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n931), .A2(new_n949), .A3(new_n942), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n672), .A2(new_n675), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT108), .B(G1981), .Z(new_n970));
  NOR2_X1   g545(.A1(G305), .A2(new_n970), .ZN(new_n971));
  OR3_X1    g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n955), .B1(new_n894), .B2(new_n936), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(G288), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT52), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n665), .B2(G1976), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n975), .B(new_n978), .C1(new_n977), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT55), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n892), .A2(KEYINPUT45), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(new_n921), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G1971), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n927), .A2(new_n894), .A3(new_n928), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G2090), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n981), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n989), .A2(new_n983), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n985), .B2(new_n711), .ZN(new_n993));
  INV_X1    g568(.A(G1961), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n987), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n711), .A2(KEYINPUT53), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n938), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G171), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n966), .A2(new_n967), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G288), .A2(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n971), .B1(new_n975), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n974), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n991), .A2(new_n981), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n956), .A2(G168), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n992), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n992), .B2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n963), .A2(new_n965), .ZN(new_n1010));
  INV_X1    g585(.A(G1956), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n987), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT110), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(KEYINPUT110), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n984), .A2(new_n921), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n985), .A2(KEYINPUT114), .A3(new_n1015), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1013), .A2(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT111), .B(KEYINPUT57), .Z(new_n1022));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n554), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n558), .B1(new_n554), .B2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1027), .B(KEYINPUT113), .C1(new_n1028), .C2(G299), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1022), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n552), .A2(new_n553), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n523), .A2(G91), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n557), .B1(new_n1034), .B2(KEYINPUT112), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1035), .B2(new_n1024), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G299), .A2(new_n1028), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1029), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1021), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n987), .A2(new_n707), .ZN(new_n1042));
  INV_X1    g617(.A(G2067), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n894), .A2(new_n936), .A3(KEYINPUT115), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n894), .A2(new_n936), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(G2067), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n589), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT116), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1039), .A2(new_n1020), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1040), .A2(new_n1041), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1039), .A2(new_n1020), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1039), .A2(new_n1020), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1048), .A2(new_n589), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1049), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n543), .A2(KEYINPUT119), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n984), .A2(new_n901), .A3(new_n921), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(KEYINPUT118), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(KEYINPUT118), .B1(new_n1046), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n589), .A2(new_n1057), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1065), .A2(KEYINPUT59), .B1(new_n1048), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1065), .A2(KEYINPUT59), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1059), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1056), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1051), .B2(KEYINPUT61), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT120), .B(new_n1053), .C1(new_n1039), .C2(new_n1020), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1052), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT54), .B1(new_n997), .B2(G171), .ZN(new_n1076));
  INV_X1    g651(.A(new_n984), .ZN(new_n1077));
  OR4_X1    g652(.A1(new_n913), .A2(new_n1077), .A3(new_n996), .A4(new_n893), .ZN(new_n1078));
  AOI21_X1  g653(.A(G301), .B1(new_n995), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT127), .B(KEYINPUT54), .Z(new_n1081));
  NAND3_X1  g656(.A1(new_n995), .A2(G301), .A3(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n998), .B2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1080), .A2(new_n992), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1075), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1009), .B1(new_n1010), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n907), .B1(new_n1000), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n896), .B(KEYINPUT48), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(new_n906), .ZN(new_n1089));
  INV_X1    g664(.A(new_n903), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n897), .B1(new_n1090), .B2(new_n752), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT46), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n897), .B2(new_n901), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n895), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(KEYINPUT47), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n785), .A2(new_n1043), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n697), .A2(new_n700), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n904), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1089), .B(new_n1096), .C1(new_n897), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1087), .A2(new_n1100), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g676(.A1(new_n847), .A2(new_n840), .ZN(new_n1103));
  NAND2_X1  g677(.A1(new_n888), .A2(new_n885), .ZN(new_n1104));
  NOR4_X1   g678(.A1(G229), .A2(new_n457), .A3(G401), .A4(G227), .ZN(new_n1105));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(G225));
  INV_X1    g680(.A(G225), .ZN(G308));
endmodule


